module notes_sequence_Mario_1(
	input clk,
	input [10:0] address,
	output reg [4:0] note,
	output reg note_on,
	output reg [12:0] delay
);

reg [18:0] note_;

always @(posedge clk) begin
case(address)
0:note_<=19'b1001110000000001010;
1:note_<=19'b0001110010000010000;
2:note_<=19'b1001110000000000001;
3:note_<=19'b0001110001111111011;
4:note_<=19'b1001110001111110101;
5:note_<=19'b0001110001111110100;
6:note_<=19'b1001110010000011100;
7:note_<=19'b0001110001111111011;
8:note_<=19'b1001110000000000001;
9:note_<=19'b0001110001111110011;
10:note_<=19'b1011001001111110110;
11:note_<=19'b0011000010000011010;
12:note_<=19'b1011000101111100110;
13:note_<=19'b0011000010000011010;
14:note_<=19'b1010010011111110001;
15:note_<=19'b0010010001111110100;
16:note_<=19'b1001010100000011000;
17:note_<=19'b0001010001111110011;
18:note_<=19'b1010100100000010001;
19:note_<=19'b0010100001111111011;
20:note_<=19'b1011000001111110101;
21:note_<=19'b0011000001111110100;
22:note_<=19'b1010110010000011100;
23:note_<=19'b0010110001111111011;
24:note_<=19'b1010100000000000001;
25:note_<=19'b0010100001111110011;
26:note_<=19'b1010010001111110110;
27:note_<=19'b0010010001011000000;
28:note_<=19'b1100010001010101011;
29:note_<=19'b0100010001010101001;
30:note_<=19'b1101010001010101100;
31:note_<=19'b0101010001010010101;
32:note_<=19'b1101100001010101011;
33:note_<=19'b0101100010000011010;
34:note_<=19'b1100110001111111101;
35:note_<=19'b0100110001111110011;
36:note_<=19'b1101010000000000001;
37:note_<=19'b0101010001111110100;
38:note_<=19'b1100010010000011100;
39:note_<=19'b0100010001111111011;
40:note_<=19'b1011100001111110101;
41:note_<=19'b0011100001111110100;
42:note_<=19'b1100000000000000001;
43:note_<=19'b0100000010000011010;
44:note_<=19'b1011000000000000001;
45:note_<=19'b0011000001111111011;
46:note_<=19'b1011000011111101010;
47:note_<=19'b0011000010000011010;
48:note_<=19'b1010010011111110001;
49:note_<=19'b0010010001111110100;
50:note_<=19'b1001010100000011000;
51:note_<=19'b0001010001111110011;
52:note_<=19'b1010100100000010001;
53:note_<=19'b0010100001111111011;
54:note_<=19'b1011000001111110101;
55:note_<=19'b0011000001111110100;
56:note_<=19'b1010110010000011100;
57:note_<=19'b0010110001111111011;
58:note_<=19'b1010100000000000001;
59:note_<=19'b0010100001111110011;
60:note_<=19'b1010010001111110110;
61:note_<=19'b0010010001011000000;
62:note_<=19'b1100010001010101011;
63:note_<=19'b0100010001010101001;
64:note_<=19'b1101010001010101100;
65:note_<=19'b0101010001010010101;
66:note_<=19'b1101100001010101011;
67:note_<=19'b0101100010000011010;
68:note_<=19'b1100110001111111101;
69:note_<=19'b0100110001111110011;
70:note_<=19'b1101010000000000001;
71:note_<=19'b0101010001111110100;
72:note_<=19'b1100010010000011100;
73:note_<=19'b0100010001111111011;
74:note_<=19'b1011100001111110101;
75:note_<=19'b0011100001111110100;
76:note_<=19'b1100000000000000001;
77:note_<=19'b0100000010000011010;
78:note_<=19'b1011000000000000001;
79:note_<=19'b0011000001111111011;
80:note_<=19'b1001010011111101010;
81:note_<=19'b0001010010000011010;
82:note_<=19'b1011000011111110001;
83:note_<=19'b0011000001111110100;
84:note_<=19'b1100010100000011000;
85:note_<=19'b0100010001111110011;
86:note_<=19'b1010100001111110110;
87:note_<=19'b0010100010000011010;
88:note_<=19'b1100010011111110001;
89:note_<=19'b0100010001111110100;
90:note_<=19'b1100010000000000001;
91:note_<=19'b0100010010000011010;
92:note_<=19'b1010100001111111101;
93:note_<=19'b0010100001111110011;
94:note_<=19'b1001010001111110110;
95:note_<=19'b0001010010000011010;
96:note_<=19'b1010010011111110001;
97:note_<=19'b0010010001111110100;
98:note_<=19'b1011000100000011000;
99:note_<=19'b0011000001111110011;
100:note_<=19'b1100010000000000001;
101:note_<=19'b0100010001111110100;
102:note_<=19'b1011001100000011000;
103:note_<=19'b0011000001111110011;
104:note_<=19'b1001010001111110110;
105:note_<=19'b0001010010000011010;
106:note_<=19'b1011000011111110001;
107:note_<=19'b0011000001111110100;
108:note_<=19'b1100010100000011000;
109:note_<=19'b0100010001111110011;
110:note_<=19'b1010100001111110110;
111:note_<=19'b0010100010000011010;
112:note_<=19'b1100010011111110001;
113:note_<=19'b0100010001111110100;
114:note_<=19'b1100010000000000001;
115:note_<=19'b0100010010000011010;
116:note_<=19'b1010100001111111101;
117:note_<=19'b0010100001111110011;
118:note_<=19'b1001010001111110110;
119:note_<=19'b0001010010000011010;
120:note_<=19'b1011010001111111101;
121:note_<=19'b0011010001111110011;
122:note_<=19'b1011110100000010001;
123:note_<=19'b0011110001111111011;
124:note_<=19'b1100010011111101010;
125:note_<=19'b0100010010000011010;
126:note_<=19'b1011000011111110001;
127:note_<=19'b0011000001111110100;
128:note_<=19'b1011000000000000001;
129:note_<=19'b0011000010000011010;
130:note_<=19'b1001010001111111101;
131:note_<=19'b0001010001111110011;
132:note_<=19'b1001010001111110110;
133:note_<=19'b0001010010000011010;
134:note_<=19'b1011000011111110001;
135:note_<=19'b0011000001111110100;
136:note_<=19'b1100010100000011000;
137:note_<=19'b0100010001111110011;
138:note_<=19'b1010100001111110110;
139:note_<=19'b0010100010000011010;
140:note_<=19'b1100010011111110001;
141:note_<=19'b0100010001111110100;
142:note_<=19'b1100010000000000001;
143:note_<=19'b0100010010000011010;
144:note_<=19'b1010100001111111101;
145:note_<=19'b0010100001111110011;
146:note_<=19'b1001010001111110110;
147:note_<=19'b0001010010000011010;
148:note_<=19'b1010010011111110001;
149:note_<=19'b0010010001111110100;
150:note_<=19'b1011000100000011000;
151:note_<=19'b0011000001111110011;
152:note_<=19'b1100010000000000001;
153:note_<=19'b0100010001111110100;
154:note_<=19'b1011001100000011000;
155:note_<=19'b0011000001111110011;
156:note_<=19'b1001010001111110110;
157:note_<=19'b0001010010000011010;
158:note_<=19'b1011000011111110001;
159:note_<=19'b0011000001111110100;
160:note_<=19'b1100010100000011000;
161:note_<=19'b0100010001111110011;
162:note_<=19'b1010100001111110110;
163:note_<=19'b0010100010000011010;
164:note_<=19'b1100010011111110001;
165:note_<=19'b0100010001111110100;
166:note_<=19'b1100010000000000001;
167:note_<=19'b0100010010000011010;
168:note_<=19'b1010100001111111101;
169:note_<=19'b0010100001111110011;
170:note_<=19'b1001010001111110110;
171:note_<=19'b0001010010000011010;
172:note_<=19'b1011010001111111101;
173:note_<=19'b0011010001111110011;
174:note_<=19'b1011110100000010001;
175:note_<=19'b0011110001111111011;
176:note_<=19'b1100010011111101010;
177:note_<=19'b0100010010000011010;
178:note_<=19'b1011000011111110001;
179:note_<=19'b0011000001111110100;
180:note_<=19'b1011000000000000001;
181:note_<=19'b0011000010000011010;
182:note_<=19'b1001010001111111101;
183:note_<=19'b0001010001111110011;
184:note_<=19'b1000010001111110110;
185:note_<=19'b0000010010000011010;
186:note_<=19'b1010000011111110001;
187:note_<=19'b0010000001111110100;
188:note_<=19'b1011010100000011000;
189:note_<=19'b0011010001111110011;
190:note_<=19'b1011000001111110110;
191:note_<=19'b0011000010000011010;
192:note_<=19'b1001010011111110001;
193:note_<=19'b0001010001111110100;
194:note_<=19'b1000000100000011000;
195:note_<=19'b0000000001111110011;
196:note_<=19'b1000010001111110110;
197:note_<=19'b0000010010000011010;
198:note_<=19'b1010000011111110001;
199:note_<=19'b0010000001111110100;
200:note_<=19'b1011010100000011000;
201:note_<=19'b0011010001111110011;
202:note_<=19'b1011000001111110110;
203:note_<=19'b0011000010000011010;
204:note_<=19'b1001010011111110001;
205:note_<=19'b0001010001111110100;
206:note_<=19'b1000000100000011000;
207:note_<=19'b0000000001111110011;
208:note_<=19'b1000010001111110110;
209:note_<=19'b0000010010000011010;
210:note_<=19'b1010000011111110001;
211:note_<=19'b0010000001111110100;
212:note_<=19'b1011010100000011000;
213:note_<=19'b0011010001111110011;
214:note_<=19'b1011000001111110110;
215:note_<=19'b0011000010000011010;
216:note_<=19'b1001010011111110001;
217:note_<=19'b0001010001111110100;
218:note_<=19'b1000000100000011000;
219:note_<=19'b0000000001111110011;
220:note_<=19'b1001110001111110110;
221:note_<=19'b0001110010000011010;
222:note_<=19'b1001110000000000001;
223:note_<=19'b0001110001111111011;
224:note_<=19'b1001110001111110101;
225:note_<=19'b0001110001111110100;
226:note_<=19'b1001110010000011100;
227:note_<=19'b0001110001111111011;
228:note_<=19'b1001110000000000001;
229:note_<=19'b0001110001111110011;
230:note_<=19'b1011001001111110110;
231:note_<=19'b0011000010000011010;
232:note_<=19'b1011000101111100110;
233:note_<=19'b0011000010000011010;
234:note_<=19'b1010010011111110001;
235:note_<=19'b0010010001111110100;
236:note_<=19'b1001010100000011000;
237:note_<=19'b0001010001111110011;
238:note_<=19'b1010100100000010001;
239:note_<=19'b0010100001111111011;
240:note_<=19'b1011000001111110101;
241:note_<=19'b0011000001111110100;
242:note_<=19'b1010110010000011100;
243:note_<=19'b0010110001111111011;
244:note_<=19'b1010100000000000001;
245:note_<=19'b0010100001111110011;
246:note_<=19'b1010010001111110110;
247:note_<=19'b0010010001011000000;
248:note_<=19'b1100010001010101011;
249:note_<=19'b0100010001010101001;
250:note_<=19'b1101010001010101100;
251:note_<=19'b0101010001010010101;
252:note_<=19'b1101100001010101011;
253:note_<=19'b0101100010000011010;
254:note_<=19'b1100110001111111101;
255:note_<=19'b0100110001111110011;
256:note_<=19'b1101010000000000001;
257:note_<=19'b0101010001111110100;
258:note_<=19'b1100010010000011100;
259:note_<=19'b0100010001111111011;
260:note_<=19'b1011100001111110101;
261:note_<=19'b0011100001111110100;
262:note_<=19'b1100000000000000001;
263:note_<=19'b0100000010000011010;
264:note_<=19'b1011000000000000001;
265:note_<=19'b0011000001111111011;
266:note_<=19'b1011000011111101010;
267:note_<=19'b0011000010000011010;
268:note_<=19'b1010010011111110001;
269:note_<=19'b0010010001111110100;
270:note_<=19'b1001010100000011000;
271:note_<=19'b0001010001111110011;
272:note_<=19'b1010100100000010001;
273:note_<=19'b0010100001111111011;
274:note_<=19'b1011000001111110101;
275:note_<=19'b0011000001111110100;
276:note_<=19'b1010110010000011100;
277:note_<=19'b0010110001111111011;
278:note_<=19'b1010100000000000001;
279:note_<=19'b0010100001111110011;
280:note_<=19'b1010010001111110110;
281:note_<=19'b0010010001011000000;
282:note_<=19'b1100010001010101011;
283:note_<=19'b0100010001010101001;
284:note_<=19'b1101010001010101100;
285:note_<=19'b0101010001010010101;
286:note_<=19'b1101100001010101011;
287:note_<=19'b0101100010000011010;
288:note_<=19'b1100110001111111101;
289:note_<=19'b0100110001111110011;
290:note_<=19'b1101010000000000001;
291:note_<=19'b0101010001111110100;
292:note_<=19'b1100010010000011100;
293:note_<=19'b0100010001111111011;
294:note_<=19'b1011100001111110101;
295:note_<=19'b0011100001111110100;
296:note_<=19'b1100000000000000001;
297:note_<=19'b0100000010000011010;
298:note_<=19'b1011000000000000001;
299:note_<=19'b0011000001111111011;
300:note_<=19'b1001010011111101010;
301:note_<=19'b0001010010000011010;
302:note_<=19'b1010110011111110001;
303:note_<=19'b0010110001111110100;
304:note_<=19'b1011000000000000001;
305:note_<=19'b0011000010000011010;
306:note_<=19'b1100010001111111101;
307:note_<=19'b0100010001111110011;
308:note_<=19'b1010100001111110110;
309:note_<=19'b0010100010000011010;
310:note_<=19'b1010100001111111101;
311:note_<=19'b0010100001111110011;
312:note_<=19'b1100010001111110110;
313:note_<=19'b0100010010000011010;
314:note_<=19'b1100010000000000001;
315:note_<=19'b0100010001111111011;
316:note_<=19'b1010100000000000001;
317:note_<=19'b0010100001111110011;
318:note_<=19'b1001110001111110110;
319:note_<=19'b0001110010000011010;
320:note_<=19'b1010100011111110001;
321:note_<=19'b0010100001111110100;
322:note_<=19'b1011000000000000001;
323:note_<=19'b0011000010000011010;
324:note_<=19'b1100000001111111101;
325:note_<=19'b0100000001111110011;
326:note_<=19'b1011000001111110110;
327:note_<=19'b0011000010000011010;
328:note_<=19'b1011000001111111101;
329:note_<=19'b0011000001111110011;
330:note_<=19'b1100010001111110110;
331:note_<=19'b0100010010000011010;
332:note_<=19'b1100010000000000001;
333:note_<=19'b0100010001111111011;
334:note_<=19'b1011000000000000001;
335:note_<=19'b0011000001111110011;
336:note_<=19'b1001010001111110110;
337:note_<=19'b0001010010000011010;
338:note_<=19'b1010110011111110001;
339:note_<=19'b0010110001111110100;
340:note_<=19'b1011000000000000001;
341:note_<=19'b0011000010000011010;
342:note_<=19'b1100010001111111101;
343:note_<=19'b0100010001111110011;
344:note_<=19'b1010100001111110110;
345:note_<=19'b0010100010000011010;
346:note_<=19'b1010100001111111101;
347:note_<=19'b0010100001111110011;
348:note_<=19'b1100010001111110110;
349:note_<=19'b0100010010000011010;
350:note_<=19'b1100010000000000001;
351:note_<=19'b0100010001111111011;
352:note_<=19'b1010100000000000001;
353:note_<=19'b0010100001111110011;
354:note_<=19'b1011000001111110110;
355:note_<=19'b0011000010000011010;
356:note_<=19'b1011000011111110001;
357:note_<=19'b0011000001111110100;
358:note_<=19'b1011000000000000001;
359:note_<=19'b0011000001011000000;
360:note_<=19'b1011100001010101011;
361:note_<=19'b0011100001010101001;
362:note_<=19'b1100000001010101100;
363:note_<=19'b0100000001010010101;
364:note_<=19'b1100010001010101011;
365:note_<=19'b0100010010000011010;
366:note_<=19'b1011000001111111101;
367:note_<=19'b0011000001111110011;
368:note_<=19'b1001010001111110110;
369:note_<=19'b0001010010000011010;
370:note_<=19'b1001010101111100110;
371:note_<=19'b0001010010000011010;
372:note_<=19'b1010110011111110001;
373:note_<=19'b0010110001111110100;
374:note_<=19'b1011000000000000001;
375:note_<=19'b0011000010000011010;
376:note_<=19'b1100010001111111101;
377:note_<=19'b0100010001111110011;
378:note_<=19'b1010100001111110110;
379:note_<=19'b0010100010000011010;
380:note_<=19'b1010100001111111101;
381:note_<=19'b0010100001111110011;
382:note_<=19'b1100010001111110110;
383:note_<=19'b0100010010000011010;
384:note_<=19'b1100010000000000001;
385:note_<=19'b0100010001111111011;
386:note_<=19'b1010100000000000001;
387:note_<=19'b0010100001111110011;
388:note_<=19'b1001110001111110110;
389:note_<=19'b0001110010000011010;
390:note_<=19'b1010100011111110001;
391:note_<=19'b0010100001111110100;
392:note_<=19'b1011000000000000001;
393:note_<=19'b0011000010000011010;
394:note_<=19'b1100000001111111101;
395:note_<=19'b0100000001111110011;
396:note_<=19'b1011000001111110110;
397:note_<=19'b0011000010000011010;
398:note_<=19'b1011000001111111101;
399:note_<=19'b0011000001111110011;
400:note_<=19'b1100010001111110110;
401:note_<=19'b0100010010000011010;
402:note_<=19'b1100010000000000001;
403:note_<=19'b0100010001111111011;
404:note_<=19'b1011000000000000001;
405:note_<=19'b0011000001111110011;
406:note_<=19'b1001010001111110110;
407:note_<=19'b0001010010000011010;
408:note_<=19'b1010110011111110001;
409:note_<=19'b0010110001111110100;
410:note_<=19'b1011000000000000001;
411:note_<=19'b0011000010000011010;
412:note_<=19'b1100010001111111101;
413:note_<=19'b0100010001111110011;
414:note_<=19'b1010100001111110110;
415:note_<=19'b0010100010000011010;
416:note_<=19'b1010100001111111101;
417:note_<=19'b0010100001111110011;
418:note_<=19'b1100010001111110110;
419:note_<=19'b0100010010000011010;
420:note_<=19'b1100010000000000001;
421:note_<=19'b0100010001111111011;
422:note_<=19'b1010100000000000001;
423:note_<=19'b0010100001111110011;
424:note_<=19'b1011000001111110110;
425:note_<=19'b0011000010000011010;
426:note_<=19'b1011000011111110001;
427:note_<=19'b0011000001111110100;
428:note_<=19'b1011000000000000001;
429:note_<=19'b0011000001011000000;
430:note_<=19'b1011100001010101011;
431:note_<=19'b0011100001010101001;
432:note_<=19'b1100000001010101100;
433:note_<=19'b0100000001010010101;
434:note_<=19'b1100010001010101011;
435:note_<=19'b0100010010000011010;
436:note_<=19'b1011000001111111101;
437:note_<=19'b0011000001111110011;
438:note_<=19'b1001010001111110110;
439:note_<=19'b0001010010000011010;
440:note_<=19'b1000010101111100110;
441:note_<=19'b0000010010000011010;
442:note_<=19'b1010000011111110001;
443:note_<=19'b0010000001111110100;
444:note_<=19'b1011010100000011000;
445:note_<=19'b0011010001111110011;
446:note_<=19'b1011000001111110110;
447:note_<=19'b0011000010000011010;
448:note_<=19'b1001010011111110001;
449:note_<=19'b0001010001111110100;
450:note_<=19'b1000000100000011000;
451:note_<=19'b0000000001111110011;
452:note_<=19'b1000010001111110110;
453:note_<=19'b0000010010000011010;
454:note_<=19'b1010000011111110001;
455:note_<=19'b0010000001111110100;
456:note_<=19'b1011010100000011000;
457:note_<=19'b0011010001111110011;
458:note_<=19'b1011000001111110110;
459:note_<=19'b0011000010000011010;
460:note_<=19'b1001010011111110001;
461:note_<=19'b0001010001111110100;
462:note_<=19'b1000000100000011000;
463:note_<=19'b0000000001111110011;
464:note_<=19'b1000010001111110110;
465:note_<=19'b0000010010000011010;
466:note_<=19'b1010000011111110001;
467:note_<=19'b0010000001111110100;
468:note_<=19'b1011010100000011000;
469:note_<=19'b0011010001111110011;
470:note_<=19'b1011000001111110110;
471:note_<=19'b0011000010000011010;
472:note_<=19'b1001010011111110001;
473:note_<=19'b0001010001111110100;
474:note_<=19'b1000000100000011000;
475:note_<=19'b0000000001111110011;
476:note_<=19'b1001110001111110110;
477:note_<=19'b0001110010000011010;
478:note_<=19'b1001110000000000001;
479:note_<=19'b0001110001111111011;
480:note_<=19'b1001110001111110101;
481:note_<=19'b0001110001111110100;
482:note_<=19'b1001110010000011100;
483:note_<=19'b0001110001111111011;
484:note_<=19'b1001110000000000001;
485:note_<=19'b0001110001111110011;
486:note_<=19'b1011001001111110110;
487:note_<=19'b0011000010000011010;
488:note_<=19'b1001010101111100110;
489:note_<=19'b0001010010000011010;
490:note_<=19'b1010110011111110001;
491:note_<=19'b0010110001111110100;
492:note_<=19'b1011000000000000001;
493:note_<=19'b0011000010000011010;
494:note_<=19'b1100010001111111101;
495:note_<=19'b0100010001111110011;
496:note_<=19'b1010100001111110110;
497:note_<=19'b0010100010000011010;
498:note_<=19'b1010100001111111101;
499:note_<=19'b0010100001111110011;
500:note_<=19'b1100010001111110110;
501:note_<=19'b0100010010000011010;
502:note_<=19'b1100010000000000001;
503:note_<=19'b0100010001111111011;
504:note_<=19'b1010100000000000001;
505:note_<=19'b0010100001111110011;
506:note_<=19'b1001110001111110110;
507:note_<=19'b0001110010000011010;
508:note_<=19'b1010100011111110001;
509:note_<=19'b0010100001111110100;
510:note_<=19'b1011000000000000001;
511:note_<=19'b0011000010000011010;
512:note_<=19'b1100000001111111101;
513:note_<=19'b0100000001111110011;
514:note_<=19'b1011000001111110110;
515:note_<=19'b0011000010000011010;
516:note_<=19'b1011000001111111101;
517:note_<=19'b0011000001111110011;
518:note_<=19'b1100010001111110110;
519:note_<=19'b0100010010000011010;
520:note_<=19'b1100010000000000001;
521:note_<=19'b0100010001111111011;
522:note_<=19'b1011000000000000001;
523:note_<=19'b0011000001111110011;
524:note_<=19'b1001010001111110110;
525:note_<=19'b0001010010000011010;
526:note_<=19'b1010110011111110001;
527:note_<=19'b0010110001111110100;
528:note_<=19'b1011000000000000001;
529:note_<=19'b0011000010000011010;
530:note_<=19'b1100010001111111101;
531:note_<=19'b0100010001111110011;
532:note_<=19'b1010100001111110110;
533:note_<=19'b0010100010000011010;
534:note_<=19'b1010100001111111101;
535:note_<=19'b0010100001111110011;
536:note_<=19'b1100010001111110110;
537:note_<=19'b0100010010000011010;
538:note_<=19'b1100010000000000001;
539:note_<=19'b0100010001111111011;
540:note_<=19'b1010100000000000001;
541:note_<=19'b0010100001111110011;
542:note_<=19'b1011000001111110110;
543:note_<=19'b0011000010000011010;
544:note_<=19'b1011000011111110001;
545:note_<=19'b0011000001111110100;
546:note_<=19'b1011000000000000001;
547:note_<=19'b0011000001011000000;
548:note_<=19'b1011100001010101011;
549:note_<=19'b0011100001010101001;
550:note_<=19'b1100000001010101100;
551:note_<=19'b0100000001010010101;
552:note_<=19'b1100010001010101011;
553:note_<=19'b0100010010000011010;
554:note_<=19'b1011000001111111101;
555:note_<=19'b0011000001111110011;
556:note_<=19'b1001010001111110110;
557:note_<=19'b0001010010000011010;
558:note_<=19'b1011000101111100110;
559:note_<=19'b0011000010000011010;
560:note_<=19'b1010010011111110001;
561:note_<=19'b0010010001111110100;
562:note_<=19'b1001010100000011000;
563:note_<=19'b0001010001111110011;
564:note_<=19'b1010100100000010001;
565:note_<=19'b0010100001111111011;
566:note_<=19'b1011000001111110101;
567:note_<=19'b0011000001111110100;
568:note_<=19'b1010110010000011100;
569:note_<=19'b0010110001111111011;
570:note_<=19'b1010100000000000001;
571:note_<=19'b0010100001111110011;
572:note_<=19'b1010010001111110110;
573:note_<=19'b0010010001011000000;
574:note_<=19'b1100010001010101011;
575:note_<=19'b0100010001010101001;
576:note_<=19'b1101010001010101100;
577:note_<=19'b0101010001010010101;
578:note_<=19'b1101100001010101011;
579:note_<=19'b0101100010000011010;
580:note_<=19'b1100110001111111101;
581:note_<=19'b0100110001111110011;
582:note_<=19'b1101010000000000001;
583:note_<=19'b0101010001111110100;
584:note_<=19'b1100010010000011100;
585:note_<=19'b0100010001111111011;
586:note_<=19'b1011100001111110101;
587:note_<=19'b0011100001111110100;
588:note_<=19'b1100000000000000001;
589:note_<=19'b0100000010000011010;
590:note_<=19'b1011000000000000001;
591:note_<=19'b0011000001111111011;
592:note_<=19'b1011000011111101010;
593:note_<=19'b0011000010000011010;
594:note_<=19'b1010010011111110001;
595:note_<=19'b0010010001111110100;
596:note_<=19'b1001010100000011000;
597:note_<=19'b0001010001111110011;
598:note_<=19'b1010100100000010001;
599:note_<=19'b0010100001111111011;
600:note_<=19'b1011000001111110101;
601:note_<=19'b0011000001111110100;
602:note_<=19'b1010110010000011100;
603:note_<=19'b0010110001111111011;
604:note_<=19'b1010100000000000001;
605:note_<=19'b0010100001111110011;
606:note_<=19'b1010010001111110110;
607:note_<=19'b0010010001011000000;
608:note_<=19'b1100010001010101011;
609:note_<=19'b0100010001010101001;
610:note_<=19'b1101010001010101100;
611:note_<=19'b0101010001010010101;
612:note_<=19'b1101100001010101011;
613:note_<=19'b0101100010000011010;
614:note_<=19'b1100110001111111101;
615:note_<=19'b0100110001111110011;
616:note_<=19'b1101010000000000001;
617:note_<=19'b0101010001111110100;
618:note_<=19'b1100010010000011100;
619:note_<=19'b0100010001111111011;
620:note_<=19'b1011100001111110101;
621:note_<=19'b0011100001111110100;
622:note_<=19'b1100000000000000001;
623:note_<=19'b0100000010000011010;
624:note_<=19'b1011000000000000001;
625:note_<=19'b0011000001111111011;
626:note_<=19'b1001010011111101010;
627:note_<=19'b0001010010000011010;
628:note_<=19'b1011000011111110001;
629:note_<=19'b0011000001111110100;
630:note_<=19'b1100010100000011000;
631:note_<=19'b0100010001111110011;
632:note_<=19'b1010100001111110110;
633:note_<=19'b0010100010000011010;
634:note_<=19'b1100010011111110001;
635:note_<=19'b0100010001111110100;
636:note_<=19'b1100010000000000001;
637:note_<=19'b0100010010000011010;
638:note_<=19'b1010100001111111101;
639:note_<=19'b0010100001111110011;
640:note_<=19'b1001010001111110110;
641:note_<=19'b0001010010000011010;
642:note_<=19'b1010010011111110001;
643:note_<=19'b0010010001111110100;
644:note_<=19'b1011000100000011000;
645:note_<=19'b0011000001111110011;
646:note_<=19'b1100010000000000001;
647:note_<=19'b0100010001111110100;
648:note_<=19'b1011001100000011000;
649:note_<=19'b0011000001111110011;
650:note_<=19'b1001010001111110110;
651:note_<=19'b0001010010000011010;
652:note_<=19'b1011000011111110001;
653:note_<=19'b0011000001111110100;
654:note_<=19'b1100010100000011000;
655:note_<=19'b0100010001111110011;
656:note_<=19'b1010100001111110110;
657:note_<=19'b0010100010000011010;
658:note_<=19'b1100010011111110001;
659:note_<=19'b0100010001111110100;
660:note_<=19'b1100010000000000001;
661:note_<=19'b0100010010000011010;
662:note_<=19'b1010100001111111101;
663:note_<=19'b0010100001111110011;
664:note_<=19'b1001010001111110110;
665:note_<=19'b0001010010000011010;
666:note_<=19'b1011010001111111101;
667:note_<=19'b0011010001111110011;
668:note_<=19'b1011110100000010001;
669:note_<=19'b0011110001111111011;
670:note_<=19'b1100010011111101010;
671:note_<=19'b0100010010000011010;
672:note_<=19'b1011000011111110001;
673:note_<=19'b0011000001111110100;
674:note_<=19'b1011000000000000001;
675:note_<=19'b0011000010000011010;
676:note_<=19'b1001010001111111101;
677:note_<=19'b0001010001111110011;
678:note_<=19'b1001010001111110110;
679:note_<=19'b0001010010000011010;
680:note_<=19'b1011000011111110001;
681:note_<=19'b0011000001111110100;
682:note_<=19'b1100010100000011000;
683:note_<=19'b0100010001111110011;
684:note_<=19'b1010100001111110110;
685:note_<=19'b0010100010000011010;
686:note_<=19'b1100010011111110001;
687:note_<=19'b0100010001111110100;
688:note_<=19'b1100010000000000001;
689:note_<=19'b0100010010000011010;
690:note_<=19'b1010100001111111101;
691:note_<=19'b0010100001111110011;
692:note_<=19'b1001010001111110110;
693:note_<=19'b0001010010000011010;
694:note_<=19'b1010010011111110001;
695:note_<=19'b0010010001111110100;
696:note_<=19'b1011000100000011000;
697:note_<=19'b0011000001111110011;
698:note_<=19'b1100010000000000001;
699:note_<=19'b0100010001111110100;
700:note_<=19'b1011001100000011000;
701:note_<=19'b0011000001111110011;
702:note_<=19'b1001010001111110110;
703:note_<=19'b0001010010000011010;
704:note_<=19'b1011000011111110001;
705:note_<=19'b0011000001111110100;
706:note_<=19'b1100010100000011000;
707:note_<=19'b0100010001111110011;
708:note_<=19'b1010100001111110110;
709:note_<=19'b0010100010000011010;
710:note_<=19'b1100010011111110001;
711:note_<=19'b0100010001111110100;
712:note_<=19'b1100010000000000001;
713:note_<=19'b0100010010000011010;
714:note_<=19'b1010100001111111101;
715:note_<=19'b0010100001111110011;
716:note_<=19'b1001010001111110110;
717:note_<=19'b0001010010000011010;
718:note_<=19'b1011010001111111101;
719:note_<=19'b0011010001111110011;
720:note_<=19'b1011110100000010001;
721:note_<=19'b0011110001111111011;
722:note_<=19'b1100010011111101010;
723:note_<=19'b0100010010000011010;
724:note_<=19'b1011000011111110001;
725:note_<=19'b0011000001111110100;
726:note_<=19'b1011000000000000001;
727:note_<=19'b0011000010000011010;
728:note_<=19'b1001010001111111101;
729:note_<=19'b0001010001111110011;
730:note_<=19'b1000010001111110110;
731:note_<=19'b0000010010000011010;
732:note_<=19'b1010000011111110001;
733:note_<=19'b0010000001111110100;
734:note_<=19'b1011010100000011000;
735:note_<=19'b0011010001111110011;
736:note_<=19'b1011000001111110110;
737:note_<=19'b0011000010000011010;
738:note_<=19'b1001010011111110001;
739:note_<=19'b0001010001111110100;
740:note_<=19'b1000000100000011000;
741:note_<=19'b0000000001111110011;
742:note_<=19'b1000010001111110110;
743:note_<=19'b0000010010000011010;
744:note_<=19'b1010000011111110001;
745:note_<=19'b0010000001111110100;
746:note_<=19'b1011010100000011000;
747:note_<=19'b0011010001111110011;
748:note_<=19'b1011000001111110110;
749:note_<=19'b0011000010000011010;
750:note_<=19'b1001010011111110001;
751:note_<=19'b0001010001111110100;
752:note_<=19'b1000000100000011000;
753:note_<=19'b0000000001111110011;
754:note_<=19'b1000010001111110110;
755:note_<=19'b0000010010000011010;
756:note_<=19'b1010000011111110001;
757:note_<=19'b0010000001111110100;
758:note_<=19'b1011010100000011000;
759:note_<=19'b0011010001111110011;
760:note_<=19'b1011000001111110110;
761:note_<=19'b0011000010000011010;
762:note_<=19'b1001010011111110001;
763:note_<=19'b0001010001111110100;
764:note_<=19'b1000000100000011000;
765:note_<=19'b0000000001111110011;
766:note_<=19'b1001110001111110110;
767:note_<=19'b0001110010000011010;
768:note_<=19'b1001110000000000001;
769:note_<=19'b0001110001111111011;
770:note_<=19'b1001110001111110101;
771:note_<=19'b0001110001111110100;
772:note_<=19'b1001110010000011100;
773:note_<=19'b0001110001111111011;
774:note_<=19'b1001110000000000001;
775:note_<=19'b0001110001111110011;
776:note_<=19'b1011001001111110110;
777:note_<=19'b0011000010000011010;
778:note_<=19'b1011000101111100110;
779:note_<=19'b0011000010000011010;
780:note_<=19'b1010010011111110001;
781:note_<=19'b0010010001111110100;
782:note_<=19'b1001010100000011000;
783:note_<=19'b0001010001111110011;
784:note_<=19'b1010100100000010001;
785:note_<=19'b0010100001111111011;
786:note_<=19'b1011000001111110101;
787:note_<=19'b0011000001111110100;
788:note_<=19'b1010110010000011100;
789:note_<=19'b0010110001111111011;
790:note_<=19'b1010100000000000001;
791:note_<=19'b0010100001111110011;
792:note_<=19'b1010010001111110110;
793:note_<=19'b0010010001011000000;
794:note_<=19'b1100010001010101011;
795:note_<=19'b0100010001010101001;
796:note_<=19'b1101010001010101100;
797:note_<=19'b0101010001010010101;
798:note_<=19'b1101100001010101011;
799:note_<=19'b0101100010000011010;
800:note_<=19'b1100110001111111101;
801:note_<=19'b0100110001111110011;
802:note_<=19'b1101010000000000001;
803:note_<=19'b0101010001111110100;
804:note_<=19'b1100010010000011100;
805:note_<=19'b0100010001111111011;
806:note_<=19'b1011100001111110101;
807:note_<=19'b0011100001111110100;
808:note_<=19'b1100000000000000001;
809:note_<=19'b0100000010000011010;
810:note_<=19'b1011000000000000001;
811:note_<=19'b0011000001111111011;
812:note_<=19'b1011000011111101010;
813:note_<=19'b0011000010000011010;
814:note_<=19'b1010010011111110001;
815:note_<=19'b0010010001111110100;
816:note_<=19'b1001010100000011000;
817:note_<=19'b0001010001111110011;
818:note_<=19'b1010100100000010001;
819:note_<=19'b0010100001111111011;
820:note_<=19'b1011000001111110101;
821:note_<=19'b0011000001111110100;
822:note_<=19'b1010110010000011100;
823:note_<=19'b0010110001111111011;
824:note_<=19'b1010100000000000001;
825:note_<=19'b0010100001111110011;
826:note_<=19'b1010010001111110110;
827:note_<=19'b0010010001011000000;
828:note_<=19'b1100010001010101011;
829:note_<=19'b0100010001010101001;
830:note_<=19'b1101010001010101100;
831:note_<=19'b0101010001010010101;
832:note_<=19'b1101100001010101011;
833:note_<=19'b0101100010000011010;
834:note_<=19'b1100110001111111101;
835:note_<=19'b0100110001111110011;
836:note_<=19'b1101010000000000001;
837:note_<=19'b0101010001111110100;
838:note_<=19'b1100010010000011100;
839:note_<=19'b0100010001111111011;
840:note_<=19'b1011100001111110101;
841:note_<=19'b0011100001111110100;
842:note_<=19'b1100000000000000001;
843:note_<=19'b0100000010000011010;
844:note_<=19'b1011000000000000001;
845:note_<=19'b0011000001111111011;
846:note_<=19'b1001010011111101010;
847:note_<=19'b0001010010000011010;
848:note_<=19'b1010110011111110001;
849:note_<=19'b0010110001111110100;
850:note_<=19'b1011000000000000001;
851:note_<=19'b0011000010000011010;
852:note_<=19'b1100010001111111101;
853:note_<=19'b0100010001111110011;
854:note_<=19'b1010100001111110110;
855:note_<=19'b0010100010000011010;
856:note_<=19'b1010100001111111101;
857:note_<=19'b0010100001111110011;
858:note_<=19'b1100010001111110110;
859:note_<=19'b0100010010000011010;
860:note_<=19'b1100010000000000001;
861:note_<=19'b0100010001111111011;
862:note_<=19'b1010100000000000001;
863:note_<=19'b0010100001111110011;
864:note_<=19'b1001110001111110110;
865:note_<=19'b0001110010000011010;
866:note_<=19'b1010100011111110001;
867:note_<=19'b0010100001111110100;
868:note_<=19'b1011000000000000001;
869:note_<=19'b0011000010000011010;
870:note_<=19'b1100000001111111101;
871:note_<=19'b0100000001111110011;
872:note_<=19'b1011000001111110110;
873:note_<=19'b0011000010000011010;
874:note_<=19'b1011000001111111101;
875:note_<=19'b0011000001111110011;
876:note_<=19'b1100010001111110110;
877:note_<=19'b0100010010000011010;
878:note_<=19'b1100010000000000001;
879:note_<=19'b0100010001111111011;
880:note_<=19'b1011000000000000001;
881:note_<=19'b0011000001111110011;
882:note_<=19'b1001010001111110110;
883:note_<=19'b0001010010000011010;
884:note_<=19'b1010110011111110001;
885:note_<=19'b0010110001111110100;
886:note_<=19'b1011000000000000001;
887:note_<=19'b0011000010000011010;
888:note_<=19'b1100010001111111101;
889:note_<=19'b0100010001111110011;
890:note_<=19'b1010100001111110110;
891:note_<=19'b0010100010000011010;
892:note_<=19'b1010100001111111101;
893:note_<=19'b0010100001111110011;
894:note_<=19'b1100010001111110110;
895:note_<=19'b0100010010000011010;
896:note_<=19'b1100010000000000001;
897:note_<=19'b0100010001111111011;
898:note_<=19'b1010100000000000001;
899:note_<=19'b0010100001111110011;
900:note_<=19'b1011000001111110110;
901:note_<=19'b0011000010000011010;
902:note_<=19'b1011000011111110001;
903:note_<=19'b0011000001111110100;
904:note_<=19'b1011000000000000001;
905:note_<=19'b0011000001011000000;
906:note_<=19'b1011100001010101011;
907:note_<=19'b0011100001010101001;
908:note_<=19'b1100000001010101100;
909:note_<=19'b0100000001010010101;
910:note_<=19'b1100010001010101011;
911:note_<=19'b0100010010000011010;
912:note_<=19'b1011000001111111101;
913:note_<=19'b0011000001111110011;
914:note_<=19'b1001010001111110110;
915:note_<=19'b0001010010000011010;
916:note_<=19'b1001010101111100110;
917:note_<=19'b0001010010000011010;
918:note_<=19'b1010110011111110001;
919:note_<=19'b0010110001111110100;
920:note_<=19'b1011000000000000001;
921:note_<=19'b0011000010000011010;
922:note_<=19'b1100010001111111101;
923:note_<=19'b0100010001111110011;
924:note_<=19'b1010100001111110110;
925:note_<=19'b0010100010000011010;
926:note_<=19'b1010100001111111101;
927:note_<=19'b0010100001111110011;
928:note_<=19'b1100010001111110110;
929:note_<=19'b0100010010000011010;
930:note_<=19'b1100010000000000001;
931:note_<=19'b0100010001111111011;
932:note_<=19'b1010100000000000001;
933:note_<=19'b0010100001111110011;
934:note_<=19'b1001110001111110110;
935:note_<=19'b0001110010000011010;
936:note_<=19'b1010100011111110001;
937:note_<=19'b0010100001111110100;
938:note_<=19'b1011000000000000001;
939:note_<=19'b0011000010000011010;
940:note_<=19'b1100000001111111101;
941:note_<=19'b0100000001111110011;
942:note_<=19'b1011000001111110110;
943:note_<=19'b0011000010000011010;
944:note_<=19'b1011000001111111101;
945:note_<=19'b0011000001111110011;
946:note_<=19'b1100010001111110110;
947:note_<=19'b0100010010000011010;
948:note_<=19'b1100010000000000001;
949:note_<=19'b0100010001111111011;
950:note_<=19'b1011000000000000001;
951:note_<=19'b0011000001111110011;
952:note_<=19'b1001010001111110110;
953:note_<=19'b0001010010000011010;
954:note_<=19'b1010110011111110001;
955:note_<=19'b0010110001111110100;
956:note_<=19'b1011000000000000001;
957:note_<=19'b0011000010000011010;
958:note_<=19'b1100010001111111101;
959:note_<=19'b0100010001111110011;
960:note_<=19'b1010100001111110110;
961:note_<=19'b0010100010000011010;
962:note_<=19'b1010100001111111101;
963:note_<=19'b0010100001111110011;
964:note_<=19'b1100010001111110110;
965:note_<=19'b0100010010000011010;
966:note_<=19'b1100010000000000001;
967:note_<=19'b0100010001111111011;
968:note_<=19'b1010100000000000001;
969:note_<=19'b0010100001111110011;
970:note_<=19'b1011000001111110110;
971:note_<=19'b0011000010000011010;
972:note_<=19'b1011000011111110001;
973:note_<=19'b0011000001111110100;
974:note_<=19'b1011000000000000001;
975:note_<=19'b0011000001011000000;
976:note_<=19'b1011100001010101011;
977:note_<=19'b0011100001010101001;
978:note_<=19'b1100000001010101100;
979:note_<=19'b0100000001010010101;
980:note_<=19'b1100010001010101011;
981:note_<=19'b0100010010000011010;
982:note_<=19'b1011000001111111101;
983:note_<=19'b0011000001111110011;
984:note_<=19'b1001010001111110110;
985:note_<=19'b0001010010000011010;
986:note_<=19'b1000010101111100110;
987:note_<=19'b0000010010000011010;
988:note_<=19'b1010000011111110001;
989:note_<=19'b0010000001111110100;
990:note_<=19'b1011010100000011000;
991:note_<=19'b0011010001111110011;
992:note_<=19'b1011000001111110110;
993:note_<=19'b0011000010000011010;
994:note_<=19'b1001010011111110001;
995:note_<=19'b0001010001111110100;
996:note_<=19'b1000000100000011000;
997:note_<=19'b0000000001111110011;
998:note_<=19'b1000010001111110110;
999:note_<=19'b0000010010000011010;
1000:note_<=19'b1010000011111110001;
1001:note_<=19'b0010000001111110100;
1002:note_<=19'b1011010100000011000;
1003:note_<=19'b0011010001111110011;
1004:note_<=19'b1011000001111110110;
1005:note_<=19'b0011000010000011010;
1006:note_<=19'b1001010011111110001;
1007:note_<=19'b0001010001111110100;
1008:note_<=19'b1000000100000011000;
1009:note_<=19'b0000000001111110011;
1010:note_<=19'b1000010001111110110;
1011:note_<=19'b0000010010000011010;
1012:note_<=19'b1010000011111110001;
1013:note_<=19'b0010000001111110100;
1014:note_<=19'b1011010100000011000;
1015:note_<=19'b0011010001111110011;
1016:note_<=19'b1011000001111110110;
1017:note_<=19'b0011000010000011010;
1018:note_<=19'b1001010011111110001;
1019:note_<=19'b0001010001111110100;
1020:note_<=19'b1000000100000011000;
1021:note_<=19'b0000000001111110011;
1022:note_<=19'b1001110001111110110;
1023:note_<=19'b0001110010000011010;
1024:note_<=19'b1001110000000000001;
1025:note_<=19'b0001110001111111011;
1026:note_<=19'b1001110001111110101;
1027:note_<=19'b0001110001111110100;
1028:note_<=19'b1001110010000011100;
1029:note_<=19'b0001110001111111011;
1030:note_<=19'b1001110000000000001;
1031:note_<=19'b0001110001111110011;
1032:note_<=19'b1011001001111110110;
1033:note_<=19'b0011000010000011010;
1034:note_<=19'b1001010101111100110;
1035:note_<=19'b0001010010000011010;
1036:note_<=19'b1010110011111110001;
1037:note_<=19'b0010110001111110100;
1038:note_<=19'b1011000000000000001;
1039:note_<=19'b0011000010000011010;
1040:note_<=19'b1100010001111111101;
1041:note_<=19'b0100010001111110011;
1042:note_<=19'b1010100001111110110;
1043:note_<=19'b0010100010000011010;
1044:note_<=19'b1010100001111111101;
1045:note_<=19'b0010100001111110011;
1046:note_<=19'b1100010001111110110;
1047:note_<=19'b0100010010000011010;
1048:note_<=19'b1100010000000000001;
1049:note_<=19'b0100010001111111011;
1050:note_<=19'b1010100000000000001;
1051:note_<=19'b0010100001111110011;
1052:note_<=19'b1001110001111110110;
1053:note_<=19'b0001110010000011010;
1054:note_<=19'b1010100011111110001;
1055:note_<=19'b0010100001111110100;
1056:note_<=19'b1011000000000000001;
1057:note_<=19'b0011000010000011010;
1058:note_<=19'b1100000001111111101;
1059:note_<=19'b0100000001111110011;
1060:note_<=19'b1011000001111110110;
1061:note_<=19'b0011000010000011010;
1062:note_<=19'b1011000001111111101;
1063:note_<=19'b0011000001111110011;
1064:note_<=19'b1100010001111110110;
1065:note_<=19'b0100010010000011010;
1066:note_<=19'b1100010000000000001;
1067:note_<=19'b0100010001111111011;
1068:note_<=19'b1011000000000000001;
1069:note_<=19'b0011000001111110011;
1070:note_<=19'b1001010001111110110;
1071:note_<=19'b0001010010000011010;
1072:note_<=19'b1010110011111110001;
1073:note_<=19'b0010110001111110100;
1074:note_<=19'b1011000000000000001;
1075:note_<=19'b0011000010000011010;
1076:note_<=19'b1100010001111111101;
1077:note_<=19'b0100010001111110011;
1078:note_<=19'b1010100001111110110;
1079:note_<=19'b0010100010000011010;
1080:note_<=19'b1010100001111111101;
1081:note_<=19'b0010100001111110011;
1082:note_<=19'b1100010001111110110;
1083:note_<=19'b0100010010000011010;
1084:note_<=19'b1100010000000000001;
1085:note_<=19'b0100010001111111011;
1086:note_<=19'b1010100000000000001;
1087:note_<=19'b0010100001111110011;
1088:note_<=19'b1011000001111110110;
1089:note_<=19'b0011000010000011010;
1090:note_<=19'b1011000011111110001;
1091:note_<=19'b0011000001111110100;
1092:note_<=19'b1011000000000000001;
1093:note_<=19'b0011000001011000000;
1094:note_<=19'b1011100001010101011;
1095:note_<=19'b0011100001010101001;
1096:note_<=19'b1100000001010101100;
1097:note_<=19'b0100000001010010101;
1098:note_<=19'b1100010001010101011;
1099:note_<=19'b0100010010000011010;
1100:note_<=19'b1011000001111111101;
1101:note_<=19'b0011000001111110011;
1102:note_<=19'b1001010001111110110;
1103:note_<=19'b0001010010000011010;
default: note_ <= 19'b0;
endcase

note_on <= note_[18:18];
note <= note_[17:13];
delay <= note_[12:0];
end
endmodule


