module notes_sequence_Mario_0(
	input clk,
	input [11:0] address,
	output reg [4:0] note,
	output reg note_on,
	output reg [13:0] delay
);

reg [19:0] note_;

always @(posedge clk) begin
case(address)
0:note_<=20'b10101100000000001010;
1:note_<=20'b11010100000000000000;
2:note_<=20'b00101100010000010000;
3:note_<=20'b01010100000000000000;
4:note_<=20'b10101100000000000001;
5:note_<=20'b11010100000000000000;
6:note_<=20'b00101100001111111011;
7:note_<=20'b01010100000000000000;
8:note_<=20'b10101100001111110101;
9:note_<=20'b11010100000000000000;
10:note_<=20'b00101100001111110100;
11:note_<=20'b01010100000000000000;
12:note_<=20'b10101100010000011100;
13:note_<=20'b11000100000000000000;
14:note_<=20'b00101100001111111011;
15:note_<=20'b01000100000000000000;
16:note_<=20'b10101100000000000001;
17:note_<=20'b11010100000000000000;
18:note_<=20'b00101100001111110011;
19:note_<=20'b01010100000000000000;
20:note_<=20'b10110000001111110110;
21:note_<=20'b11000000000000000000;
22:note_<=20'b11100000000000000000;
23:note_<=20'b00110000010000011010;
24:note_<=20'b01000000000000000000;
25:note_<=20'b01100000000000000000;
26:note_<=20'b10110000101111100110;
27:note_<=20'b00110000010000011010;
28:note_<=20'b10100100101111100110;
29:note_<=20'b11000100000000000000;
30:note_<=20'b00100100010000011010;
31:note_<=20'b01000100000000000000;
32:note_<=20'b10010100011111110001;
33:note_<=20'b10110000000000000000;
34:note_<=20'b00010100001111110100;
35:note_<=20'b00110000000000000000;
36:note_<=20'b10000000100000011000;
37:note_<=20'b10100100000000000000;
38:note_<=20'b00000000001111110011;
39:note_<=20'b00100100000000000000;
40:note_<=20'b10010100100000010001;
41:note_<=20'b10111000000000000000;
42:note_<=20'b00010100001111111011;
43:note_<=20'b00111000000000000000;
44:note_<=20'b10011100001111110101;
45:note_<=20'b11000000000000000000;
46:note_<=20'b00011100001111110100;
47:note_<=20'b01000000000000000000;
48:note_<=20'b10011000010000011100;
49:note_<=20'b10111100000000000000;
50:note_<=20'b00011000001111111011;
51:note_<=20'b00111100000000000000;
52:note_<=20'b10010100000000000001;
53:note_<=20'b10111000000000000000;
54:note_<=20'b00010100001111110011;
55:note_<=20'b00111000000000000000;
56:note_<=20'b10010100001111110110;
57:note_<=20'b10110000000000000000;
58:note_<=20'b00010100001011000000;
59:note_<=20'b00110000000000000000;
60:note_<=20'b10110000001010101011;
61:note_<=20'b11010100000000000000;
62:note_<=20'b00110000001010101001;
63:note_<=20'b01010100000000000000;
64:note_<=20'b11000000001010101100;
65:note_<=20'b11100000000000000000;
66:note_<=20'b01000000001010010101;
67:note_<=20'b01100000000000000000;
68:note_<=20'b11000100001010101011;
69:note_<=20'b11101000000000000000;
70:note_<=20'b01000100010000011010;
71:note_<=20'b01101000000000000000;
72:note_<=20'b10111000001111111101;
73:note_<=20'b11011000000000000000;
74:note_<=20'b00111000001111110011;
75:note_<=20'b01011000000000000000;
76:note_<=20'b11000000000000000001;
77:note_<=20'b11100000000000000000;
78:note_<=20'b01000000001111110100;
79:note_<=20'b01100000000000000000;
80:note_<=20'b10111000010000011100;
81:note_<=20'b11010100000000000000;
82:note_<=20'b00111000001111111011;
83:note_<=20'b01010100000000000000;
84:note_<=20'b10100100001111110101;
85:note_<=20'b11000100000000000000;
86:note_<=20'b00100100001111110100;
87:note_<=20'b01000100000000000000;
88:note_<=20'b10101000000000000001;
89:note_<=20'b11001100000000000000;
90:note_<=20'b00101000010000011010;
91:note_<=20'b01001100000000000000;
92:note_<=20'b10011100000000000001;
93:note_<=20'b11000000000000000000;
94:note_<=20'b00011100001111111011;
95:note_<=20'b01000000000000000000;
96:note_<=20'b10100100011111101010;
97:note_<=20'b11000100000000000000;
98:note_<=20'b00100100010000011010;
99:note_<=20'b01000100000000000000;
100:note_<=20'b10010100011111110001;
101:note_<=20'b10110000000000000000;
102:note_<=20'b00010100001111110100;
103:note_<=20'b00110000000000000000;
104:note_<=20'b10000000100000011000;
105:note_<=20'b10100100000000000000;
106:note_<=20'b00000000001111110011;
107:note_<=20'b00100100000000000000;
108:note_<=20'b10010100100000010001;
109:note_<=20'b10111000000000000000;
110:note_<=20'b00010100001111111011;
111:note_<=20'b00111000000000000000;
112:note_<=20'b10011100001111110101;
113:note_<=20'b11000000000000000000;
114:note_<=20'b00011100001111110100;
115:note_<=20'b01000000000000000000;
116:note_<=20'b10011000010000011100;
117:note_<=20'b10111100000000000000;
118:note_<=20'b00011000001111111011;
119:note_<=20'b00111100000000000000;
120:note_<=20'b10010100000000000001;
121:note_<=20'b10111000000000000000;
122:note_<=20'b00010100001111110011;
123:note_<=20'b00111000000000000000;
124:note_<=20'b10010100001111110110;
125:note_<=20'b10110000000000000000;
126:note_<=20'b00010100001011000000;
127:note_<=20'b00110000000000000000;
128:note_<=20'b10110000001010101011;
129:note_<=20'b11010100000000000000;
130:note_<=20'b00110000001010101001;
131:note_<=20'b01010100000000000000;
132:note_<=20'b11000000001010101100;
133:note_<=20'b11100000000000000000;
134:note_<=20'b01000000001010010101;
135:note_<=20'b01100000000000000000;
136:note_<=20'b11000100001010101011;
137:note_<=20'b11101000000000000000;
138:note_<=20'b01000100010000011010;
139:note_<=20'b01101000000000000000;
140:note_<=20'b10111000001111111101;
141:note_<=20'b11011000000000000000;
142:note_<=20'b00111000001111110011;
143:note_<=20'b01011000000000000000;
144:note_<=20'b11000000000000000001;
145:note_<=20'b11100000000000000000;
146:note_<=20'b01000000001111110100;
147:note_<=20'b01100000000000000000;
148:note_<=20'b10111000010000011100;
149:note_<=20'b11010100000000000000;
150:note_<=20'b00111000001111111011;
151:note_<=20'b01010100000000000000;
152:note_<=20'b10100100001111110101;
153:note_<=20'b11000100000000000000;
154:note_<=20'b00100100001111110100;
155:note_<=20'b01000100000000000000;
156:note_<=20'b10101000000000000001;
157:note_<=20'b11001100000000000000;
158:note_<=20'b00101000010000011010;
159:note_<=20'b01001100000000000000;
160:note_<=20'b10011100000000000001;
161:note_<=20'b11000000000000000000;
162:note_<=20'b00011100001111111011;
163:note_<=20'b01000000000000000000;
164:note_<=20'b11010101000000000001;
165:note_<=20'b11100000000000000000;
166:note_<=20'b01010100001111110011;
167:note_<=20'b01100000000000000000;
168:note_<=20'b11010000000000000001;
169:note_<=20'b11011100000000000000;
170:note_<=20'b01010000001111110100;
171:note_<=20'b01011100000000000000;
172:note_<=20'b11001100000000000001;
173:note_<=20'b11011000000000000000;
174:note_<=20'b01001100010000011010;
175:note_<=20'b01011000000000000000;
176:note_<=20'b11000000000000000001;
177:note_<=20'b11010000000000000000;
178:note_<=20'b01000000001111111011;
179:note_<=20'b01010000000000000000;
180:note_<=20'b11000100001111110101;
181:note_<=20'b11010100000000000000;
182:note_<=20'b01000100001111110100;
183:note_<=20'b01010100000000000000;
184:note_<=20'b10100100010000011100;
185:note_<=20'b10110100000000000000;
186:note_<=20'b00100100001111111011;
187:note_<=20'b00110100000000000000;
188:note_<=20'b10101000000000000001;
189:note_<=20'b10111000000000000000;
190:note_<=20'b00101000001111110011;
191:note_<=20'b00111000000000000000;
192:note_<=20'b10110000000000000001;
193:note_<=20'b11000100000000000000;
194:note_<=20'b00110000001111110100;
195:note_<=20'b01000100000000000000;
196:note_<=20'b10010100010000011100;
197:note_<=20'b10111000000000000000;
198:note_<=20'b00010100001111111011;
199:note_<=20'b00111000000000000000;
200:note_<=20'b10100100000000000001;
201:note_<=20'b11000100000000000000;
202:note_<=20'b00100100001111110011;
203:note_<=20'b01000100000000000000;
204:note_<=20'b10101000000000000001;
205:note_<=20'b11001100000000000000;
206:note_<=20'b00101000001111110100;
207:note_<=20'b01001100000000000000;
208:note_<=20'b11010100100000011000;
209:note_<=20'b11100000000000000000;
210:note_<=20'b01010100001111110011;
211:note_<=20'b01100000000000000000;
212:note_<=20'b11010000000000000001;
213:note_<=20'b11011100000000000000;
214:note_<=20'b01010000001111110100;
215:note_<=20'b01011100000000000000;
216:note_<=20'b11001100000000000001;
217:note_<=20'b11011000000000000000;
218:note_<=20'b01001100010000011010;
219:note_<=20'b01011000000000000000;
220:note_<=20'b11000000000000000001;
221:note_<=20'b11010000000000000000;
222:note_<=20'b01000000001111111011;
223:note_<=20'b01010000000000000000;
224:note_<=20'b11000100001111110101;
225:note_<=20'b11010100000000000000;
226:note_<=20'b01000100001111110100;
227:note_<=20'b01010100000000000000;
228:note_<=20'b11011000010000011100;
229:note_<=20'b11100000000000000000;
230:note_<=20'b11110100000000000000;
231:note_<=20'b01011000001111111011;
232:note_<=20'b01100000000000000000;
233:note_<=20'b01110100000000000000;
234:note_<=20'b11011000001111110101;
235:note_<=20'b11100000000000000000;
236:note_<=20'b11110100000000000000;
237:note_<=20'b01011000001111110100;
238:note_<=20'b01100000000000000000;
239:note_<=20'b01110100000000000000;
240:note_<=20'b11011000000000000001;
241:note_<=20'b11100000000000000000;
242:note_<=20'b11110100000000000000;
243:note_<=20'b01011000010000011010;
244:note_<=20'b01100000000000000000;
245:note_<=20'b01110100000000000000;
246:note_<=20'b11010101001111111101;
247:note_<=20'b11100000000000000000;
248:note_<=20'b01010100001111110011;
249:note_<=20'b01100000000000000000;
250:note_<=20'b11010000000000000001;
251:note_<=20'b11011100000000000000;
252:note_<=20'b01010000001111110100;
253:note_<=20'b01011100000000000000;
254:note_<=20'b11001100000000000001;
255:note_<=20'b11011000000000000000;
256:note_<=20'b01001100010000011010;
257:note_<=20'b01011000000000000000;
258:note_<=20'b11000000000000000001;
259:note_<=20'b11010000000000000000;
260:note_<=20'b01000000001111111011;
261:note_<=20'b01010000000000000000;
262:note_<=20'b11000100001111110101;
263:note_<=20'b11010100000000000000;
264:note_<=20'b01000100001111110100;
265:note_<=20'b01010100000000000000;
266:note_<=20'b10100100010000011100;
267:note_<=20'b10110100000000000000;
268:note_<=20'b00100100001111111011;
269:note_<=20'b00110100000000000000;
270:note_<=20'b10101000000000000001;
271:note_<=20'b10111000000000000000;
272:note_<=20'b00101000001111110011;
273:note_<=20'b00111000000000000000;
274:note_<=20'b10110000000000000001;
275:note_<=20'b11000100000000000000;
276:note_<=20'b00110000001111110100;
277:note_<=20'b01000100000000000000;
278:note_<=20'b10010100010000011100;
279:note_<=20'b10111000000000000000;
280:note_<=20'b00010100001111111011;
281:note_<=20'b00111000000000000000;
282:note_<=20'b10100100000000000001;
283:note_<=20'b11000100000000000000;
284:note_<=20'b00100100001111110011;
285:note_<=20'b01000100000000000000;
286:note_<=20'b10101000000000000001;
287:note_<=20'b11001100000000000000;
288:note_<=20'b00101000001111110100;
289:note_<=20'b01001100000000000000;
290:note_<=20'b10110100100000011000;
291:note_<=20'b11010000000000000000;
292:note_<=20'b00110100001111110011;
293:note_<=20'b01010000000000000000;
294:note_<=20'b10101000100000010001;
295:note_<=20'b11001100000000000000;
296:note_<=20'b00101000001111111011;
297:note_<=20'b01001100000000000000;
298:note_<=20'b10100100011111101010;
299:note_<=20'b11000100000000000000;
300:note_<=20'b00100100010000011010;
301:note_<=20'b01000100000000000000;
302:note_<=20'b11010110001111111101;
303:note_<=20'b11100000000000000000;
304:note_<=20'b01010100001111110011;
305:note_<=20'b01100000000000000000;
306:note_<=20'b11010000000000000001;
307:note_<=20'b11011100000000000000;
308:note_<=20'b01010000001111110100;
309:note_<=20'b01011100000000000000;
310:note_<=20'b11001100000000000001;
311:note_<=20'b11011000000000000000;
312:note_<=20'b01001100010000011010;
313:note_<=20'b01011000000000000000;
314:note_<=20'b11000000000000000001;
315:note_<=20'b11010000000000000000;
316:note_<=20'b01000000001111111011;
317:note_<=20'b01010000000000000000;
318:note_<=20'b11000100001111110101;
319:note_<=20'b11010100000000000000;
320:note_<=20'b01000100001111110100;
321:note_<=20'b01010100000000000000;
322:note_<=20'b10100100010000011100;
323:note_<=20'b10110100000000000000;
324:note_<=20'b00100100001111111011;
325:note_<=20'b00110100000000000000;
326:note_<=20'b10101000000000000001;
327:note_<=20'b10111000000000000000;
328:note_<=20'b00101000001111110011;
329:note_<=20'b00111000000000000000;
330:note_<=20'b10110000000000000001;
331:note_<=20'b11000100000000000000;
332:note_<=20'b00110000001111110100;
333:note_<=20'b01000100000000000000;
334:note_<=20'b10010100010000011100;
335:note_<=20'b10111000000000000000;
336:note_<=20'b00010100001111111011;
337:note_<=20'b00111000000000000000;
338:note_<=20'b10100100000000000001;
339:note_<=20'b11000100000000000000;
340:note_<=20'b00100100001111110011;
341:note_<=20'b01000100000000000000;
342:note_<=20'b10101000000000000001;
343:note_<=20'b11001100000000000000;
344:note_<=20'b00101000001111110100;
345:note_<=20'b01001100000000000000;
346:note_<=20'b11010100100000011000;
347:note_<=20'b11100000000000000000;
348:note_<=20'b01010100001111110011;
349:note_<=20'b01100000000000000000;
350:note_<=20'b11010000000000000001;
351:note_<=20'b11011100000000000000;
352:note_<=20'b01010000001111110100;
353:note_<=20'b01011100000000000000;
354:note_<=20'b11001100000000000001;
355:note_<=20'b11011000000000000000;
356:note_<=20'b01001100010000011010;
357:note_<=20'b01011000000000000000;
358:note_<=20'b11000000000000000001;
359:note_<=20'b11010000000000000000;
360:note_<=20'b01000000001111111011;
361:note_<=20'b01010000000000000000;
362:note_<=20'b11000100001111110101;
363:note_<=20'b11010100000000000000;
364:note_<=20'b01000100001111110100;
365:note_<=20'b01010100000000000000;
366:note_<=20'b11011000010000011100;
367:note_<=20'b11100000000000000000;
368:note_<=20'b11110100000000000000;
369:note_<=20'b01011000001111111011;
370:note_<=20'b01100000000000000000;
371:note_<=20'b01110100000000000000;
372:note_<=20'b11011000001111110101;
373:note_<=20'b11100000000000000000;
374:note_<=20'b11110100000000000000;
375:note_<=20'b01011000001111110100;
376:note_<=20'b01100000000000000000;
377:note_<=20'b01110100000000000000;
378:note_<=20'b11011000000000000001;
379:note_<=20'b11100000000000000000;
380:note_<=20'b11110100000000000000;
381:note_<=20'b01011000010000011010;
382:note_<=20'b01100000000000000000;
383:note_<=20'b01110100000000000000;
384:note_<=20'b11010101001111111101;
385:note_<=20'b11100000000000000000;
386:note_<=20'b01010100001111110011;
387:note_<=20'b01100000000000000000;
388:note_<=20'b11010000000000000001;
389:note_<=20'b11011100000000000000;
390:note_<=20'b01010000001111110100;
391:note_<=20'b01011100000000000000;
392:note_<=20'b11001100000000000001;
393:note_<=20'b11011000000000000000;
394:note_<=20'b01001100010000011010;
395:note_<=20'b01011000000000000000;
396:note_<=20'b11000000000000000001;
397:note_<=20'b11010000000000000000;
398:note_<=20'b01000000001111111011;
399:note_<=20'b01010000000000000000;
400:note_<=20'b11000100001111110101;
401:note_<=20'b11010100000000000000;
402:note_<=20'b01000100001111110100;
403:note_<=20'b01010100000000000000;
404:note_<=20'b10100100010000011100;
405:note_<=20'b10110100000000000000;
406:note_<=20'b00100100001111111011;
407:note_<=20'b00110100000000000000;
408:note_<=20'b10101000000000000001;
409:note_<=20'b10111000000000000000;
410:note_<=20'b00101000001111110011;
411:note_<=20'b00111000000000000000;
412:note_<=20'b10110000000000000001;
413:note_<=20'b11000100000000000000;
414:note_<=20'b00110000001111110100;
415:note_<=20'b01000100000000000000;
416:note_<=20'b10010100010000011100;
417:note_<=20'b10111000000000000000;
418:note_<=20'b00010100001111111011;
419:note_<=20'b00111000000000000000;
420:note_<=20'b10100100000000000001;
421:note_<=20'b11000100000000000000;
422:note_<=20'b00100100001111110011;
423:note_<=20'b01000100000000000000;
424:note_<=20'b10101000000000000001;
425:note_<=20'b11001100000000000000;
426:note_<=20'b00101000001111110100;
427:note_<=20'b01001100000000000000;
428:note_<=20'b10110100100000011000;
429:note_<=20'b11010000000000000000;
430:note_<=20'b00110100001111110011;
431:note_<=20'b01010000000000000000;
432:note_<=20'b10101000100000010001;
433:note_<=20'b11001100000000000000;
434:note_<=20'b00101000001111111011;
435:note_<=20'b01001100000000000000;
436:note_<=20'b10100100011111101010;
437:note_<=20'b11000100000000000000;
438:note_<=20'b00100100010000011010;
439:note_<=20'b01000100000000000000;
440:note_<=20'b10110101101111100110;
441:note_<=20'b11000100000000000000;
442:note_<=20'b00110100010000011010;
443:note_<=20'b01000100000000000000;
444:note_<=20'b10110100000000000001;
445:note_<=20'b11000100000000000000;
446:note_<=20'b00110100001111111011;
447:note_<=20'b01000100000000000000;
448:note_<=20'b10110100001111110101;
449:note_<=20'b11000100000000000000;
450:note_<=20'b00110100001111110100;
451:note_<=20'b01000100000000000000;
452:note_<=20'b10110100010000011100;
453:note_<=20'b11000100000000000000;
454:note_<=20'b00110100001111111011;
455:note_<=20'b01000100000000000000;
456:note_<=20'b10111100000000000001;
457:note_<=20'b11001100000000000000;
458:note_<=20'b00111100001111110011;
459:note_<=20'b01001100000000000000;
460:note_<=20'b10110000001111110110;
461:note_<=20'b11010100000000000000;
462:note_<=20'b00110000010000011010;
463:note_<=20'b01010100000000000000;
464:note_<=20'b10100100000000000001;
465:note_<=20'b11000100000000000000;
466:note_<=20'b00100100001111111011;
467:note_<=20'b01000100000000000000;
468:note_<=20'b10100100001111110101;
469:note_<=20'b10111000000000000000;
470:note_<=20'b00100100001111110100;
471:note_<=20'b00111000000000000000;
472:note_<=20'b10010100000000000001;
473:note_<=20'b10110000000000000000;
474:note_<=20'b00010100010000011010;
475:note_<=20'b00110000000000000000;
476:note_<=20'b10110100101111100110;
477:note_<=20'b11000100000000000000;
478:note_<=20'b00110100010000011010;
479:note_<=20'b01000100000000000000;
480:note_<=20'b10110100000000000001;
481:note_<=20'b11000100000000000000;
482:note_<=20'b00110100001111111011;
483:note_<=20'b01000100000000000000;
484:note_<=20'b10110100001111110101;
485:note_<=20'b11000100000000000000;
486:note_<=20'b00110100001111110100;
487:note_<=20'b01000100000000000000;
488:note_<=20'b10110100010000011100;
489:note_<=20'b11000100000000000000;
490:note_<=20'b00110100001111111011;
491:note_<=20'b01000100000000000000;
492:note_<=20'b10111100000000000001;
493:note_<=20'b11001100000000000000;
494:note_<=20'b00111100001111110011;
495:note_<=20'b01001100000000000000;
496:note_<=20'b10110000000000000001;
497:note_<=20'b11010100000000000000;
498:note_<=20'b00110000001111110100;
499:note_<=20'b01010100000000000000;
500:note_<=20'b10110110000000000001;
501:note_<=20'b11000100000000000000;
502:note_<=20'b00110100010000011010;
503:note_<=20'b01000100000000000000;
504:note_<=20'b10110100000000000001;
505:note_<=20'b11000100000000000000;
506:note_<=20'b00110100001111111011;
507:note_<=20'b01000100000000000000;
508:note_<=20'b10110100001111110101;
509:note_<=20'b11000100000000000000;
510:note_<=20'b00110100001111110100;
511:note_<=20'b01000100000000000000;
512:note_<=20'b10110100010000011100;
513:note_<=20'b11000100000000000000;
514:note_<=20'b00110100001111111011;
515:note_<=20'b01000100000000000000;
516:note_<=20'b10111100000000000001;
517:note_<=20'b11001100000000000000;
518:note_<=20'b00111100001111110011;
519:note_<=20'b01001100000000000000;
520:note_<=20'b10110000001111110110;
521:note_<=20'b11010100000000000000;
522:note_<=20'b00110000010000011010;
523:note_<=20'b01010100000000000000;
524:note_<=20'b10100100000000000001;
525:note_<=20'b11000100000000000000;
526:note_<=20'b00100100001111111011;
527:note_<=20'b01000100000000000000;
528:note_<=20'b10100100001111110101;
529:note_<=20'b10111000000000000000;
530:note_<=20'b00100100001111110100;
531:note_<=20'b00111000000000000000;
532:note_<=20'b10010100000000000001;
533:note_<=20'b10110000000000000000;
534:note_<=20'b00010100010000011010;
535:note_<=20'b00110000000000000000;
536:note_<=20'b10101100101111100110;
537:note_<=20'b11010100000000000000;
538:note_<=20'b00101100010000011010;
539:note_<=20'b01010100000000000000;
540:note_<=20'b10101100000000000001;
541:note_<=20'b11010100000000000000;
542:note_<=20'b00101100001111111011;
543:note_<=20'b01010100000000000000;
544:note_<=20'b10101100001111110101;
545:note_<=20'b11010100000000000000;
546:note_<=20'b00101100001111110100;
547:note_<=20'b01010100000000000000;
548:note_<=20'b10101100010000011100;
549:note_<=20'b11000100000000000000;
550:note_<=20'b00101100001111111011;
551:note_<=20'b01000100000000000000;
552:note_<=20'b10101100000000000001;
553:note_<=20'b11010100000000000000;
554:note_<=20'b00101100001111110011;
555:note_<=20'b01010100000000000000;
556:note_<=20'b10110000001111110110;
557:note_<=20'b11000000000000000000;
558:note_<=20'b11100000000000000000;
559:note_<=20'b00110000010000011010;
560:note_<=20'b01000000000000000000;
561:note_<=20'b01100000000000000000;
562:note_<=20'b10110000101111100110;
563:note_<=20'b00110000010000011010;
564:note_<=20'b10100100101111100110;
565:note_<=20'b11000100000000000000;
566:note_<=20'b00100100010000011010;
567:note_<=20'b01000100000000000000;
568:note_<=20'b10010100011111110001;
569:note_<=20'b10110000000000000000;
570:note_<=20'b00010100001111110100;
571:note_<=20'b00110000000000000000;
572:note_<=20'b10000000100000011000;
573:note_<=20'b10100100000000000000;
574:note_<=20'b00000000001111110011;
575:note_<=20'b00100100000000000000;
576:note_<=20'b10010100100000010001;
577:note_<=20'b10111000000000000000;
578:note_<=20'b00010100001111111011;
579:note_<=20'b00111000000000000000;
580:note_<=20'b10011100001111110101;
581:note_<=20'b11000000000000000000;
582:note_<=20'b00011100001111110100;
583:note_<=20'b01000000000000000000;
584:note_<=20'b10011000010000011100;
585:note_<=20'b10111100000000000000;
586:note_<=20'b00011000001111111011;
587:note_<=20'b00111100000000000000;
588:note_<=20'b10010100000000000001;
589:note_<=20'b10111000000000000000;
590:note_<=20'b00010100001111110011;
591:note_<=20'b00111000000000000000;
592:note_<=20'b10010100001111110110;
593:note_<=20'b10110000000000000000;
594:note_<=20'b00010100001011000000;
595:note_<=20'b00110000000000000000;
596:note_<=20'b10110000001010101011;
597:note_<=20'b11010100000000000000;
598:note_<=20'b00110000001010101001;
599:note_<=20'b01010100000000000000;
600:note_<=20'b11000000001010101100;
601:note_<=20'b11100000000000000000;
602:note_<=20'b01000000001010010101;
603:note_<=20'b01100000000000000000;
604:note_<=20'b11000100001010101011;
605:note_<=20'b11101000000000000000;
606:note_<=20'b01000100010000011010;
607:note_<=20'b01101000000000000000;
608:note_<=20'b10111000001111111101;
609:note_<=20'b11011000000000000000;
610:note_<=20'b00111000001111110011;
611:note_<=20'b01011000000000000000;
612:note_<=20'b11000000000000000001;
613:note_<=20'b11100000000000000000;
614:note_<=20'b01000000001111110100;
615:note_<=20'b01100000000000000000;
616:note_<=20'b10111000010000011100;
617:note_<=20'b11010100000000000000;
618:note_<=20'b00111000001111111011;
619:note_<=20'b01010100000000000000;
620:note_<=20'b10100100001111110101;
621:note_<=20'b11000100000000000000;
622:note_<=20'b00100100001111110100;
623:note_<=20'b01000100000000000000;
624:note_<=20'b10101000000000000001;
625:note_<=20'b11001100000000000000;
626:note_<=20'b00101000010000011010;
627:note_<=20'b01001100000000000000;
628:note_<=20'b10011100000000000001;
629:note_<=20'b11000000000000000000;
630:note_<=20'b00011100001111111011;
631:note_<=20'b01000000000000000000;
632:note_<=20'b10100100011111101010;
633:note_<=20'b11000100000000000000;
634:note_<=20'b00100100010000011010;
635:note_<=20'b01000100000000000000;
636:note_<=20'b10010100011111110001;
637:note_<=20'b10110000000000000000;
638:note_<=20'b00010100001111110100;
639:note_<=20'b00110000000000000000;
640:note_<=20'b10000000100000011000;
641:note_<=20'b10100100000000000000;
642:note_<=20'b00000000001111110011;
643:note_<=20'b00100100000000000000;
644:note_<=20'b10010100100000010001;
645:note_<=20'b10111000000000000000;
646:note_<=20'b00010100001111111011;
647:note_<=20'b00111000000000000000;
648:note_<=20'b10011100001111110101;
649:note_<=20'b11000000000000000000;
650:note_<=20'b00011100001111110100;
651:note_<=20'b01000000000000000000;
652:note_<=20'b10011000010000011100;
653:note_<=20'b10111100000000000000;
654:note_<=20'b00011000001111111011;
655:note_<=20'b00111100000000000000;
656:note_<=20'b10010100000000000001;
657:note_<=20'b10111000000000000000;
658:note_<=20'b00010100001111110011;
659:note_<=20'b00111000000000000000;
660:note_<=20'b10010100001111110110;
661:note_<=20'b10110000000000000000;
662:note_<=20'b00010100001011000000;
663:note_<=20'b00110000000000000000;
664:note_<=20'b10110000001010101011;
665:note_<=20'b11010100000000000000;
666:note_<=20'b00110000001010101001;
667:note_<=20'b01010100000000000000;
668:note_<=20'b11000000001010101100;
669:note_<=20'b11100000000000000000;
670:note_<=20'b01000000001010010101;
671:note_<=20'b01100000000000000000;
672:note_<=20'b11000100001010101011;
673:note_<=20'b11101000000000000000;
674:note_<=20'b01000100010000011010;
675:note_<=20'b01101000000000000000;
676:note_<=20'b10111000001111111101;
677:note_<=20'b11011000000000000000;
678:note_<=20'b00111000001111110011;
679:note_<=20'b01011000000000000000;
680:note_<=20'b11000000000000000001;
681:note_<=20'b11100000000000000000;
682:note_<=20'b01000000001111110100;
683:note_<=20'b01100000000000000000;
684:note_<=20'b10111000010000011100;
685:note_<=20'b11010100000000000000;
686:note_<=20'b00111000001111111011;
687:note_<=20'b01010100000000000000;
688:note_<=20'b10100100001111110101;
689:note_<=20'b11000100000000000000;
690:note_<=20'b00100100001111110100;
691:note_<=20'b01000100000000000000;
692:note_<=20'b10101000000000000001;
693:note_<=20'b11001100000000000000;
694:note_<=20'b00101000010000011010;
695:note_<=20'b01001100000000000000;
696:note_<=20'b10011100000000000001;
697:note_<=20'b11000000000000000000;
698:note_<=20'b00011100001111111011;
699:note_<=20'b01000000000000000000;
700:note_<=20'b11000100011111101010;
701:note_<=20'b11010100000000000000;
702:note_<=20'b01000100010000011010;
703:note_<=20'b01010100000000000000;
704:note_<=20'b10111000000000000001;
705:note_<=20'b11000100000000000000;
706:note_<=20'b00111000001111111011;
707:note_<=20'b01000100000000000000;
708:note_<=20'b10100100001111110101;
709:note_<=20'b10110000000000000000;
710:note_<=20'b00100100001111110100;
711:note_<=20'b00110000000000000000;
712:note_<=20'b10100100100000011000;
713:note_<=20'b10110100000000000000;
714:note_<=20'b00100100001111110011;
715:note_<=20'b00110100000000000000;
716:note_<=20'b10101000001111110110;
717:note_<=20'b10111000000000000000;
718:note_<=20'b00101000010000011010;
719:note_<=20'b00111000000000000000;
720:note_<=20'b11000100000000000001;
721:note_<=20'b11011000000000000000;
722:note_<=20'b01000100001111111011;
723:note_<=20'b01011000000000000000;
724:note_<=20'b11000100001111110101;
725:note_<=20'b11011000000000000000;
726:note_<=20'b01000100001111110100;
727:note_<=20'b01011000000000000000;
728:note_<=20'b10101000000000000001;
729:note_<=20'b10111000000000000000;
730:note_<=20'b00101000010000011010;
731:note_<=20'b00111000000000000000;
732:note_<=20'b10110000101111100110;
733:note_<=20'b11000000000000000000;
734:note_<=20'b00110000001011000000;
735:note_<=20'b01000000000000000000;
736:note_<=20'b11011000001010101011;
737:note_<=20'b11101000000000000000;
738:note_<=20'b01011000001010101001;
739:note_<=20'b01101000000000000000;
740:note_<=20'b11011000001010101100;
741:note_<=20'b11101000000000000000;
742:note_<=20'b01011000001010010101;
743:note_<=20'b01101000000000000000;
744:note_<=20'b11011000001010101011;
745:note_<=20'b11101000000000000000;
746:note_<=20'b01011000001011000000;
747:note_<=20'b01101000000000000000;
748:note_<=20'b11010100001010101011;
749:note_<=20'b11100000000000000000;
750:note_<=20'b01010100001010101001;
751:note_<=20'b01100000000000000000;
752:note_<=20'b11001100001010101100;
753:note_<=20'b11011000000000000000;
754:note_<=20'b01001100001010010101;
755:note_<=20'b01011000000000000000;
756:note_<=20'b11000100001010101011;
757:note_<=20'b11010100000000000000;
758:note_<=20'b01000100010000011010;
759:note_<=20'b01010100000000000000;
760:note_<=20'b10111000000000000001;
761:note_<=20'b11000100000000000000;
762:note_<=20'b00111000001111111011;
763:note_<=20'b01000100000000000000;
764:note_<=20'b10101000001111110101;
765:note_<=20'b10111000000000000000;
766:note_<=20'b00101000001111110100;
767:note_<=20'b00111000000000000000;
768:note_<=20'b10100100000000000001;
769:note_<=20'b10110000000000000000;
770:note_<=20'b00100100010000011010;
771:note_<=20'b00110000000000000000;
772:note_<=20'b11000100101111100110;
773:note_<=20'b11010100000000000000;
774:note_<=20'b01000100010000011010;
775:note_<=20'b01010100000000000000;
776:note_<=20'b10111000000000000001;
777:note_<=20'b11000100000000000000;
778:note_<=20'b00111000001111111011;
779:note_<=20'b01000100000000000000;
780:note_<=20'b10100100001111110101;
781:note_<=20'b10110000000000000000;
782:note_<=20'b00100100001111110100;
783:note_<=20'b00110000000000000000;
784:note_<=20'b10100100100000011000;
785:note_<=20'b10110100000000000000;
786:note_<=20'b00100100001111110011;
787:note_<=20'b00110100000000000000;
788:note_<=20'b10101000001111110110;
789:note_<=20'b10111000000000000000;
790:note_<=20'b00101000010000011010;
791:note_<=20'b00111000000000000000;
792:note_<=20'b11000100000000000001;
793:note_<=20'b11011000000000000000;
794:note_<=20'b01000100001111111011;
795:note_<=20'b01011000000000000000;
796:note_<=20'b11000100001111110101;
797:note_<=20'b11011000000000000000;
798:note_<=20'b01000100001111110100;
799:note_<=20'b01011000000000000000;
800:note_<=20'b10101000000000000001;
801:note_<=20'b10111000000000000000;
802:note_<=20'b00101000010000011010;
803:note_<=20'b00111000000000000000;
804:note_<=20'b10110000101111100110;
805:note_<=20'b11000000000000000000;
806:note_<=20'b00110000010000011010;
807:note_<=20'b01000000000000000000;
808:note_<=20'b11001100000000000001;
809:note_<=20'b11011000000000000000;
810:note_<=20'b01001100001111111011;
811:note_<=20'b01011000000000000000;
812:note_<=20'b11001100001111110101;
813:note_<=20'b11011000000000000000;
814:note_<=20'b01001100001111110100;
815:note_<=20'b01011000000000000000;
816:note_<=20'b11001100000000000001;
817:note_<=20'b11011000000000000000;
818:note_<=20'b01001100001011000000;
819:note_<=20'b01011000000000000000;
820:note_<=20'b11000100001010101011;
821:note_<=20'b11010100000000000000;
822:note_<=20'b01000100001010101001;
823:note_<=20'b01010100000000000000;
824:note_<=20'b11000000001010101100;
825:note_<=20'b11001100000000000000;
826:note_<=20'b01000000001010010101;
827:note_<=20'b01001100000000000000;
828:note_<=20'b10110000001010101011;
829:note_<=20'b11000100000000000000;
830:note_<=20'b00110000010000011010;
831:note_<=20'b01000100000000000000;
832:note_<=20'b10100100000000000001;
833:note_<=20'b00100100001111111011;
834:note_<=20'b10100100001111110101;
835:note_<=20'b00100100001111110100;
836:note_<=20'b10010100000000000001;
837:note_<=20'b00010100010000011010;
838:note_<=20'b11000100101111100110;
839:note_<=20'b11010100000000000000;
840:note_<=20'b01000100010000011010;
841:note_<=20'b01010100000000000000;
842:note_<=20'b10111000000000000001;
843:note_<=20'b11000100000000000000;
844:note_<=20'b00111000001111111011;
845:note_<=20'b01000100000000000000;
846:note_<=20'b10100100001111110101;
847:note_<=20'b10110000000000000000;
848:note_<=20'b00100100001111110100;
849:note_<=20'b00110000000000000000;
850:note_<=20'b10100100100000011000;
851:note_<=20'b10110100000000000000;
852:note_<=20'b00100100001111110011;
853:note_<=20'b00110100000000000000;
854:note_<=20'b10101000001111110110;
855:note_<=20'b10111000000000000000;
856:note_<=20'b00101000010000011010;
857:note_<=20'b00111000000000000000;
858:note_<=20'b11000100000000000001;
859:note_<=20'b11011000000000000000;
860:note_<=20'b01000100001111111011;
861:note_<=20'b01011000000000000000;
862:note_<=20'b11000100001111110101;
863:note_<=20'b11011000000000000000;
864:note_<=20'b01000100001111110100;
865:note_<=20'b01011000000000000000;
866:note_<=20'b10101000000000000001;
867:note_<=20'b10111000000000000000;
868:note_<=20'b00101000010000011010;
869:note_<=20'b00111000000000000000;
870:note_<=20'b10110000101111100110;
871:note_<=20'b11000000000000000000;
872:note_<=20'b00110000001011000000;
873:note_<=20'b01000000000000000000;
874:note_<=20'b11011000001010101011;
875:note_<=20'b11101000000000000000;
876:note_<=20'b01011000001010101001;
877:note_<=20'b01101000000000000000;
878:note_<=20'b11011000001010101100;
879:note_<=20'b11101000000000000000;
880:note_<=20'b01011000001010010101;
881:note_<=20'b01101000000000000000;
882:note_<=20'b11011000001010101011;
883:note_<=20'b11101000000000000000;
884:note_<=20'b01011000001011000000;
885:note_<=20'b01101000000000000000;
886:note_<=20'b11010100001010101011;
887:note_<=20'b11100000000000000000;
888:note_<=20'b01010100001010101001;
889:note_<=20'b01100000000000000000;
890:note_<=20'b11001100001010101100;
891:note_<=20'b11011000000000000000;
892:note_<=20'b01001100001010010101;
893:note_<=20'b01011000000000000000;
894:note_<=20'b11000100001010101011;
895:note_<=20'b11010100000000000000;
896:note_<=20'b01000100010000011010;
897:note_<=20'b01010100000000000000;
898:note_<=20'b10111000000000000001;
899:note_<=20'b11000100000000000000;
900:note_<=20'b00111000001111111011;
901:note_<=20'b01000100000000000000;
902:note_<=20'b10101000001111110101;
903:note_<=20'b10111000000000000000;
904:note_<=20'b00101000001111110100;
905:note_<=20'b00111000000000000000;
906:note_<=20'b10100100000000000001;
907:note_<=20'b10110000000000000000;
908:note_<=20'b00100100010000011010;
909:note_<=20'b00110000000000000000;
910:note_<=20'b11000100101111100110;
911:note_<=20'b11010100000000000000;
912:note_<=20'b01000100010000011010;
913:note_<=20'b01010100000000000000;
914:note_<=20'b10111000000000000001;
915:note_<=20'b11000100000000000000;
916:note_<=20'b00111000001111111011;
917:note_<=20'b01000100000000000000;
918:note_<=20'b10100100001111110101;
919:note_<=20'b10110000000000000000;
920:note_<=20'b00100100001111110100;
921:note_<=20'b00110000000000000000;
922:note_<=20'b10100100100000011000;
923:note_<=20'b10110100000000000000;
924:note_<=20'b00100100001111110011;
925:note_<=20'b00110100000000000000;
926:note_<=20'b10101000001111110110;
927:note_<=20'b10111000000000000000;
928:note_<=20'b00101000010000011010;
929:note_<=20'b00111000000000000000;
930:note_<=20'b11000100000000000001;
931:note_<=20'b11011000000000000000;
932:note_<=20'b01000100001111111011;
933:note_<=20'b01011000000000000000;
934:note_<=20'b11000100001111110101;
935:note_<=20'b11011000000000000000;
936:note_<=20'b01000100001111110100;
937:note_<=20'b01011000000000000000;
938:note_<=20'b10101000000000000001;
939:note_<=20'b10111000000000000000;
940:note_<=20'b00101000010000011010;
941:note_<=20'b00111000000000000000;
942:note_<=20'b10110000101111100110;
943:note_<=20'b11000000000000000000;
944:note_<=20'b00110000010000011010;
945:note_<=20'b01000000000000000000;
946:note_<=20'b11001100000000000001;
947:note_<=20'b11011000000000000000;
948:note_<=20'b01001100001111111011;
949:note_<=20'b01011000000000000000;
950:note_<=20'b11001100001111110101;
951:note_<=20'b11011000000000000000;
952:note_<=20'b01001100001111110100;
953:note_<=20'b01011000000000000000;
954:note_<=20'b11001100000000000001;
955:note_<=20'b11011000000000000000;
956:note_<=20'b01001100001011000000;
957:note_<=20'b01011000000000000000;
958:note_<=20'b11000100001010101011;
959:note_<=20'b11010100000000000000;
960:note_<=20'b01000100001010101001;
961:note_<=20'b01010100000000000000;
962:note_<=20'b11000000001010101100;
963:note_<=20'b11001100000000000000;
964:note_<=20'b01000000001010010101;
965:note_<=20'b01001100000000000000;
966:note_<=20'b10110000001010101011;
967:note_<=20'b11000100000000000000;
968:note_<=20'b00110000010000011010;
969:note_<=20'b01000100000000000000;
970:note_<=20'b10100100000000000001;
971:note_<=20'b00100100001111111011;
972:note_<=20'b10100100001111110101;
973:note_<=20'b00100100001111110100;
974:note_<=20'b10010100000000000001;
975:note_<=20'b00010100010000011010;
976:note_<=20'b10110100101111100110;
977:note_<=20'b11000100000000000000;
978:note_<=20'b00110100010000011010;
979:note_<=20'b01000100000000000000;
980:note_<=20'b10110100000000000001;
981:note_<=20'b11000100000000000000;
982:note_<=20'b00110100001111111011;
983:note_<=20'b01000100000000000000;
984:note_<=20'b10110100001111110101;
985:note_<=20'b11000100000000000000;
986:note_<=20'b00110100001111110100;
987:note_<=20'b01000100000000000000;
988:note_<=20'b10110100010000011100;
989:note_<=20'b11000100000000000000;
990:note_<=20'b00110100001111111011;
991:note_<=20'b01000100000000000000;
992:note_<=20'b10111100000000000001;
993:note_<=20'b11001100000000000000;
994:note_<=20'b00111100001111110011;
995:note_<=20'b01001100000000000000;
996:note_<=20'b10110000001111110110;
997:note_<=20'b11010100000000000000;
998:note_<=20'b00110000010000011010;
999:note_<=20'b01010100000000000000;
1000:note_<=20'b10100100000000000001;
1001:note_<=20'b11000100000000000000;
1002:note_<=20'b00100100001111111011;
1003:note_<=20'b01000100000000000000;
1004:note_<=20'b10100100001111110101;
1005:note_<=20'b10111000000000000000;
1006:note_<=20'b00100100001111110100;
1007:note_<=20'b00111000000000000000;
1008:note_<=20'b10010100000000000001;
1009:note_<=20'b10110000000000000000;
1010:note_<=20'b00010100010000011010;
1011:note_<=20'b00110000000000000000;
1012:note_<=20'b10110100101111100110;
1013:note_<=20'b11000100000000000000;
1014:note_<=20'b00110100010000011010;
1015:note_<=20'b01000100000000000000;
1016:note_<=20'b10110100000000000001;
1017:note_<=20'b11000100000000000000;
1018:note_<=20'b00110100001111111011;
1019:note_<=20'b01000100000000000000;
1020:note_<=20'b10110100001111110101;
1021:note_<=20'b11000100000000000000;
1022:note_<=20'b00110100001111110100;
1023:note_<=20'b01000100000000000000;
1024:note_<=20'b10110100010000011100;
1025:note_<=20'b11000100000000000000;
1026:note_<=20'b00110100001111111011;
1027:note_<=20'b01000100000000000000;
1028:note_<=20'b10111100000000000001;
1029:note_<=20'b11001100000000000000;
1030:note_<=20'b00111100001111110011;
1031:note_<=20'b01001100000000000000;
1032:note_<=20'b10110000000000000001;
1033:note_<=20'b11010100000000000000;
1034:note_<=20'b00110000001111110100;
1035:note_<=20'b01010100000000000000;
1036:note_<=20'b10110110000000000001;
1037:note_<=20'b11000100000000000000;
1038:note_<=20'b00110100010000011010;
1039:note_<=20'b01000100000000000000;
1040:note_<=20'b10110100000000000001;
1041:note_<=20'b11000100000000000000;
1042:note_<=20'b00110100001111111011;
1043:note_<=20'b01000100000000000000;
1044:note_<=20'b10110100001111110101;
1045:note_<=20'b11000100000000000000;
1046:note_<=20'b00110100001111110100;
1047:note_<=20'b01000100000000000000;
1048:note_<=20'b10110100010000011100;
1049:note_<=20'b11000100000000000000;
1050:note_<=20'b00110100001111111011;
1051:note_<=20'b01000100000000000000;
1052:note_<=20'b10111100000000000001;
1053:note_<=20'b11001100000000000000;
1054:note_<=20'b00111100001111110011;
1055:note_<=20'b01001100000000000000;
1056:note_<=20'b10110000001111110110;
1057:note_<=20'b11010100000000000000;
1058:note_<=20'b00110000010000011010;
1059:note_<=20'b01010100000000000000;
1060:note_<=20'b10100100000000000001;
1061:note_<=20'b11000100000000000000;
1062:note_<=20'b00100100001111111011;
1063:note_<=20'b01000100000000000000;
1064:note_<=20'b10100100001111110101;
1065:note_<=20'b10111000000000000000;
1066:note_<=20'b00100100001111110100;
1067:note_<=20'b00111000000000000000;
1068:note_<=20'b10010100000000000001;
1069:note_<=20'b10110000000000000000;
1070:note_<=20'b00010100010000011010;
1071:note_<=20'b00110000000000000000;
1072:note_<=20'b10101100101111100110;
1073:note_<=20'b11010100000000000000;
1074:note_<=20'b00101100010000011010;
1075:note_<=20'b01010100000000000000;
1076:note_<=20'b10101100000000000001;
1077:note_<=20'b11010100000000000000;
1078:note_<=20'b00101100001111111011;
1079:note_<=20'b01010100000000000000;
1080:note_<=20'b10101100001111110101;
1081:note_<=20'b11010100000000000000;
1082:note_<=20'b00101100001111110100;
1083:note_<=20'b01010100000000000000;
1084:note_<=20'b10101100010000011100;
1085:note_<=20'b11000100000000000000;
1086:note_<=20'b00101100001111111011;
1087:note_<=20'b01000100000000000000;
1088:note_<=20'b10101100000000000001;
1089:note_<=20'b11010100000000000000;
1090:note_<=20'b00101100001111110011;
1091:note_<=20'b01010100000000000000;
1092:note_<=20'b10110000001111110110;
1093:note_<=20'b11000000000000000000;
1094:note_<=20'b11100000000000000000;
1095:note_<=20'b00110000010000011010;
1096:note_<=20'b01000000000000000000;
1097:note_<=20'b01100000000000000000;
1098:note_<=20'b10110000101111100110;
1099:note_<=20'b00110000010000011010;
1100:note_<=20'b11000100101111100110;
1101:note_<=20'b11010100000000000000;
1102:note_<=20'b01000100010000011010;
1103:note_<=20'b01010100000000000000;
1104:note_<=20'b10111000000000000001;
1105:note_<=20'b11000100000000000000;
1106:note_<=20'b00111000001111111011;
1107:note_<=20'b01000100000000000000;
1108:note_<=20'b10100100001111110101;
1109:note_<=20'b10110000000000000000;
1110:note_<=20'b00100100001111110100;
1111:note_<=20'b00110000000000000000;
1112:note_<=20'b10100100100000011000;
1113:note_<=20'b10110100000000000000;
1114:note_<=20'b00100100001111110011;
1115:note_<=20'b00110100000000000000;
1116:note_<=20'b10101000001111110110;
1117:note_<=20'b10111000000000000000;
1118:note_<=20'b00101000010000011010;
1119:note_<=20'b00111000000000000000;
1120:note_<=20'b11000100000000000001;
1121:note_<=20'b11011000000000000000;
1122:note_<=20'b01000100001111111011;
1123:note_<=20'b01011000000000000000;
1124:note_<=20'b11000100001111110101;
1125:note_<=20'b11011000000000000000;
1126:note_<=20'b01000100001111110100;
1127:note_<=20'b01011000000000000000;
1128:note_<=20'b10101000000000000001;
1129:note_<=20'b10111000000000000000;
1130:note_<=20'b00101000010000011010;
1131:note_<=20'b00111000000000000000;
1132:note_<=20'b10110000101111100110;
1133:note_<=20'b11000000000000000000;
1134:note_<=20'b00110000001011000000;
1135:note_<=20'b01000000000000000000;
1136:note_<=20'b11011000001010101011;
1137:note_<=20'b11101000000000000000;
1138:note_<=20'b01011000001010101001;
1139:note_<=20'b01101000000000000000;
1140:note_<=20'b11011000001010101100;
1141:note_<=20'b11101000000000000000;
1142:note_<=20'b01011000001010010101;
1143:note_<=20'b01101000000000000000;
1144:note_<=20'b11011000001010101011;
1145:note_<=20'b11101000000000000000;
1146:note_<=20'b01011000001011000000;
1147:note_<=20'b01101000000000000000;
1148:note_<=20'b11010100001010101011;
1149:note_<=20'b11100000000000000000;
1150:note_<=20'b01010100001010101001;
1151:note_<=20'b01100000000000000000;
1152:note_<=20'b11001100001010101100;
1153:note_<=20'b11011000000000000000;
1154:note_<=20'b01001100001010010101;
1155:note_<=20'b01011000000000000000;
1156:note_<=20'b11000100001010101011;
1157:note_<=20'b11010100000000000000;
1158:note_<=20'b01000100010000011010;
1159:note_<=20'b01010100000000000000;
1160:note_<=20'b10111000000000000001;
1161:note_<=20'b11000100000000000000;
1162:note_<=20'b00111000001111111011;
1163:note_<=20'b01000100000000000000;
1164:note_<=20'b10101000001111110101;
1165:note_<=20'b10111000000000000000;
1166:note_<=20'b00101000001111110100;
1167:note_<=20'b00111000000000000000;
1168:note_<=20'b10100100000000000001;
1169:note_<=20'b10110000000000000000;
1170:note_<=20'b00100100010000011010;
1171:note_<=20'b00110000000000000000;
1172:note_<=20'b11000100101111100110;
1173:note_<=20'b11010100000000000000;
1174:note_<=20'b01000100010000011010;
1175:note_<=20'b01010100000000000000;
1176:note_<=20'b10111000000000000001;
1177:note_<=20'b11000100000000000000;
1178:note_<=20'b00111000001111111011;
1179:note_<=20'b01000100000000000000;
1180:note_<=20'b10100100001111110101;
1181:note_<=20'b10110000000000000000;
1182:note_<=20'b00100100001111110100;
1183:note_<=20'b00110000000000000000;
1184:note_<=20'b10100100100000011000;
1185:note_<=20'b10110100000000000000;
1186:note_<=20'b00100100001111110011;
1187:note_<=20'b00110100000000000000;
1188:note_<=20'b10101000001111110110;
1189:note_<=20'b10111000000000000000;
1190:note_<=20'b00101000010000011010;
1191:note_<=20'b00111000000000000000;
1192:note_<=20'b11000100000000000001;
1193:note_<=20'b11011000000000000000;
1194:note_<=20'b01000100001111111011;
1195:note_<=20'b01011000000000000000;
1196:note_<=20'b11000100001111110101;
1197:note_<=20'b11011000000000000000;
1198:note_<=20'b01000100001111110100;
1199:note_<=20'b01011000000000000000;
1200:note_<=20'b10101000000000000001;
1201:note_<=20'b10111000000000000000;
1202:note_<=20'b00101000010000011010;
1203:note_<=20'b00111000000000000000;
1204:note_<=20'b10110000101111100110;
1205:note_<=20'b11000000000000000000;
1206:note_<=20'b00110000010000011010;
1207:note_<=20'b01000000000000000000;
1208:note_<=20'b11001100000000000001;
1209:note_<=20'b11011000000000000000;
1210:note_<=20'b01001100001111111011;
1211:note_<=20'b01011000000000000000;
1212:note_<=20'b11001100001111110101;
1213:note_<=20'b11011000000000000000;
1214:note_<=20'b01001100001111110100;
1215:note_<=20'b01011000000000000000;
1216:note_<=20'b11001100000000000001;
1217:note_<=20'b11011000000000000000;
1218:note_<=20'b01001100001011000000;
1219:note_<=20'b01011000000000000000;
1220:note_<=20'b11000100001010101011;
1221:note_<=20'b11010100000000000000;
1222:note_<=20'b01000100001010101001;
1223:note_<=20'b01010100000000000000;
1224:note_<=20'b11000000001010101100;
1225:note_<=20'b11001100000000000000;
1226:note_<=20'b01000000001010010101;
1227:note_<=20'b01001100000000000000;
1228:note_<=20'b10110000001010101011;
1229:note_<=20'b11000100000000000000;
1230:note_<=20'b00110000010000011010;
1231:note_<=20'b01000100000000000000;
1232:note_<=20'b10100100000000000001;
1233:note_<=20'b00100100001111111011;
1234:note_<=20'b10100100001111110101;
1235:note_<=20'b00100100001111110100;
1236:note_<=20'b10010100000000000001;
1237:note_<=20'b00010100010000011010;
1238:note_<=20'b10100100101111100110;
1239:note_<=20'b11000100000000000000;
1240:note_<=20'b00100100010000011010;
1241:note_<=20'b01000100000000000000;
1242:note_<=20'b10010100011111110001;
1243:note_<=20'b10110000000000000000;
1244:note_<=20'b00010100001111110100;
1245:note_<=20'b00110000000000000000;
1246:note_<=20'b10000000100000011000;
1247:note_<=20'b10100100000000000000;
1248:note_<=20'b00000000001111110011;
1249:note_<=20'b00100100000000000000;
1250:note_<=20'b10010100100000010001;
1251:note_<=20'b10111000000000000000;
1252:note_<=20'b00010100001111111011;
1253:note_<=20'b00111000000000000000;
1254:note_<=20'b10011100001111110101;
1255:note_<=20'b11000000000000000000;
1256:note_<=20'b00011100001111110100;
1257:note_<=20'b01000000000000000000;
1258:note_<=20'b10011000010000011100;
1259:note_<=20'b10111100000000000000;
1260:note_<=20'b00011000001111111011;
1261:note_<=20'b00111100000000000000;
1262:note_<=20'b10010100000000000001;
1263:note_<=20'b10111000000000000000;
1264:note_<=20'b00010100001111110011;
1265:note_<=20'b00111000000000000000;
1266:note_<=20'b10010100001111110110;
1267:note_<=20'b10110000000000000000;
1268:note_<=20'b00010100001011000000;
1269:note_<=20'b00110000000000000000;
1270:note_<=20'b10110000001010101011;
1271:note_<=20'b11010100000000000000;
1272:note_<=20'b00110000001010101001;
1273:note_<=20'b01010100000000000000;
1274:note_<=20'b11000000001010101100;
1275:note_<=20'b11100000000000000000;
1276:note_<=20'b01000000001010010101;
1277:note_<=20'b01100000000000000000;
1278:note_<=20'b11000100001010101011;
1279:note_<=20'b11101000000000000000;
1280:note_<=20'b01000100010000011010;
1281:note_<=20'b01101000000000000000;
1282:note_<=20'b10111000001111111101;
1283:note_<=20'b11011000000000000000;
1284:note_<=20'b00111000001111110011;
1285:note_<=20'b01011000000000000000;
1286:note_<=20'b11000000000000000001;
1287:note_<=20'b11100000000000000000;
1288:note_<=20'b01000000001111110100;
1289:note_<=20'b01100000000000000000;
1290:note_<=20'b10111000010000011100;
1291:note_<=20'b11010100000000000000;
1292:note_<=20'b00111000001111111011;
1293:note_<=20'b01010100000000000000;
1294:note_<=20'b10100100001111110101;
1295:note_<=20'b11000100000000000000;
1296:note_<=20'b00100100001111110100;
1297:note_<=20'b01000100000000000000;
1298:note_<=20'b10101000000000000001;
1299:note_<=20'b11001100000000000000;
1300:note_<=20'b00101000010000011010;
1301:note_<=20'b01001100000000000000;
1302:note_<=20'b10011100000000000001;
1303:note_<=20'b11000000000000000000;
1304:note_<=20'b00011100001111111011;
1305:note_<=20'b01000000000000000000;
1306:note_<=20'b10100100011111101010;
1307:note_<=20'b11000100000000000000;
1308:note_<=20'b00100100010000011010;
1309:note_<=20'b01000100000000000000;
1310:note_<=20'b10010100011111110001;
1311:note_<=20'b10110000000000000000;
1312:note_<=20'b00010100001111110100;
1313:note_<=20'b00110000000000000000;
1314:note_<=20'b10000000100000011000;
1315:note_<=20'b10100100000000000000;
1316:note_<=20'b00000000001111110011;
1317:note_<=20'b00100100000000000000;
1318:note_<=20'b10010100100000010001;
1319:note_<=20'b10111000000000000000;
1320:note_<=20'b00010100001111111011;
1321:note_<=20'b00111000000000000000;
1322:note_<=20'b10011100001111110101;
1323:note_<=20'b11000000000000000000;
1324:note_<=20'b00011100001111110100;
1325:note_<=20'b01000000000000000000;
1326:note_<=20'b10011000010000011100;
1327:note_<=20'b10111100000000000000;
1328:note_<=20'b00011000001111111011;
1329:note_<=20'b00111100000000000000;
1330:note_<=20'b10010100000000000001;
1331:note_<=20'b10111000000000000000;
1332:note_<=20'b00010100001111110011;
1333:note_<=20'b00111000000000000000;
1334:note_<=20'b10010100001111110110;
1335:note_<=20'b10110000000000000000;
1336:note_<=20'b00010100001011000000;
1337:note_<=20'b00110000000000000000;
1338:note_<=20'b10110000001010101011;
1339:note_<=20'b11010100000000000000;
1340:note_<=20'b00110000001010101001;
1341:note_<=20'b01010100000000000000;
1342:note_<=20'b11000000001010101100;
1343:note_<=20'b11100000000000000000;
1344:note_<=20'b01000000001010010101;
1345:note_<=20'b01100000000000000000;
1346:note_<=20'b11000100001010101011;
1347:note_<=20'b11101000000000000000;
1348:note_<=20'b01000100010000011010;
1349:note_<=20'b01101000000000000000;
1350:note_<=20'b10111000001111111101;
1351:note_<=20'b11011000000000000000;
1352:note_<=20'b00111000001111110011;
1353:note_<=20'b01011000000000000000;
1354:note_<=20'b11000000000000000001;
1355:note_<=20'b11100000000000000000;
1356:note_<=20'b01000000001111110100;
1357:note_<=20'b01100000000000000000;
1358:note_<=20'b10111000010000011100;
1359:note_<=20'b11010100000000000000;
1360:note_<=20'b00111000001111111011;
1361:note_<=20'b01010100000000000000;
1362:note_<=20'b10100100001111110101;
1363:note_<=20'b11000100000000000000;
1364:note_<=20'b00100100001111110100;
1365:note_<=20'b01000100000000000000;
1366:note_<=20'b10101000000000000001;
1367:note_<=20'b11001100000000000000;
1368:note_<=20'b00101000010000011010;
1369:note_<=20'b01001100000000000000;
1370:note_<=20'b10011100000000000001;
1371:note_<=20'b11000000000000000000;
1372:note_<=20'b00011100001111111011;
1373:note_<=20'b01000000000000000000;
1374:note_<=20'b11010101000000000001;
1375:note_<=20'b11100000000000000000;
1376:note_<=20'b01010100001111110011;
1377:note_<=20'b01100000000000000000;
1378:note_<=20'b11010000000000000001;
1379:note_<=20'b11011100000000000000;
1380:note_<=20'b01010000001111110100;
1381:note_<=20'b01011100000000000000;
1382:note_<=20'b11001100000000000001;
1383:note_<=20'b11011000000000000000;
1384:note_<=20'b01001100010000011010;
1385:note_<=20'b01011000000000000000;
1386:note_<=20'b11000000000000000001;
1387:note_<=20'b11010000000000000000;
1388:note_<=20'b01000000001111111011;
1389:note_<=20'b01010000000000000000;
1390:note_<=20'b11000100001111110101;
1391:note_<=20'b11010100000000000000;
1392:note_<=20'b01000100001111110100;
1393:note_<=20'b01010100000000000000;
1394:note_<=20'b10100100010000011100;
1395:note_<=20'b10110100000000000000;
1396:note_<=20'b00100100001111111011;
1397:note_<=20'b00110100000000000000;
1398:note_<=20'b10101000000000000001;
1399:note_<=20'b10111000000000000000;
1400:note_<=20'b00101000001111110011;
1401:note_<=20'b00111000000000000000;
1402:note_<=20'b10110000000000000001;
1403:note_<=20'b11000100000000000000;
1404:note_<=20'b00110000001111110100;
1405:note_<=20'b01000100000000000000;
1406:note_<=20'b10010100010000011100;
1407:note_<=20'b10111000000000000000;
1408:note_<=20'b00010100001111111011;
1409:note_<=20'b00111000000000000000;
1410:note_<=20'b10100100000000000001;
1411:note_<=20'b11000100000000000000;
1412:note_<=20'b00100100001111110011;
1413:note_<=20'b01000100000000000000;
1414:note_<=20'b10101000000000000001;
1415:note_<=20'b11001100000000000000;
1416:note_<=20'b00101000001111110100;
1417:note_<=20'b01001100000000000000;
1418:note_<=20'b11010100100000011000;
1419:note_<=20'b11100000000000000000;
1420:note_<=20'b01010100001111110011;
1421:note_<=20'b01100000000000000000;
1422:note_<=20'b11010000000000000001;
1423:note_<=20'b11011100000000000000;
1424:note_<=20'b01010000001111110100;
1425:note_<=20'b01011100000000000000;
1426:note_<=20'b11001100000000000001;
1427:note_<=20'b11011000000000000000;
1428:note_<=20'b01001100010000011010;
1429:note_<=20'b01011000000000000000;
1430:note_<=20'b11000000000000000001;
1431:note_<=20'b11010000000000000000;
1432:note_<=20'b01000000001111111011;
1433:note_<=20'b01010000000000000000;
1434:note_<=20'b11000100001111110101;
1435:note_<=20'b11010100000000000000;
1436:note_<=20'b01000100001111110100;
1437:note_<=20'b01010100000000000000;
1438:note_<=20'b11011000010000011100;
1439:note_<=20'b11100000000000000000;
1440:note_<=20'b11110100000000000000;
1441:note_<=20'b01011000001111111011;
1442:note_<=20'b01100000000000000000;
1443:note_<=20'b01110100000000000000;
1444:note_<=20'b11011000001111110101;
1445:note_<=20'b11100000000000000000;
1446:note_<=20'b11110100000000000000;
1447:note_<=20'b01011000001111110100;
1448:note_<=20'b01100000000000000000;
1449:note_<=20'b01110100000000000000;
1450:note_<=20'b11011000000000000001;
1451:note_<=20'b11100000000000000000;
1452:note_<=20'b11110100000000000000;
1453:note_<=20'b01011000010000011010;
1454:note_<=20'b01100000000000000000;
1455:note_<=20'b01110100000000000000;
1456:note_<=20'b11010101001111111101;
1457:note_<=20'b11100000000000000000;
1458:note_<=20'b01010100001111110011;
1459:note_<=20'b01100000000000000000;
1460:note_<=20'b11010000000000000001;
1461:note_<=20'b11011100000000000000;
1462:note_<=20'b01010000001111110100;
1463:note_<=20'b01011100000000000000;
1464:note_<=20'b11001100000000000001;
1465:note_<=20'b11011000000000000000;
1466:note_<=20'b01001100010000011010;
1467:note_<=20'b01011000000000000000;
1468:note_<=20'b11000000000000000001;
1469:note_<=20'b11010000000000000000;
1470:note_<=20'b01000000001111111011;
1471:note_<=20'b01010000000000000000;
1472:note_<=20'b11000100001111110101;
1473:note_<=20'b11010100000000000000;
1474:note_<=20'b01000100001111110100;
1475:note_<=20'b01010100000000000000;
1476:note_<=20'b10100100010000011100;
1477:note_<=20'b10110100000000000000;
1478:note_<=20'b00100100001111111011;
1479:note_<=20'b00110100000000000000;
1480:note_<=20'b10101000000000000001;
1481:note_<=20'b10111000000000000000;
1482:note_<=20'b00101000001111110011;
1483:note_<=20'b00111000000000000000;
1484:note_<=20'b10110000000000000001;
1485:note_<=20'b11000100000000000000;
1486:note_<=20'b00110000001111110100;
1487:note_<=20'b01000100000000000000;
1488:note_<=20'b10010100010000011100;
1489:note_<=20'b10111000000000000000;
1490:note_<=20'b00010100001111111011;
1491:note_<=20'b00111000000000000000;
1492:note_<=20'b10100100000000000001;
1493:note_<=20'b11000100000000000000;
1494:note_<=20'b00100100001111110011;
1495:note_<=20'b01000100000000000000;
1496:note_<=20'b10101000000000000001;
1497:note_<=20'b11001100000000000000;
1498:note_<=20'b00101000001111110100;
1499:note_<=20'b01001100000000000000;
1500:note_<=20'b10110100100000011000;
1501:note_<=20'b11010000000000000000;
1502:note_<=20'b00110100001111110011;
1503:note_<=20'b01010000000000000000;
1504:note_<=20'b10101000100000010001;
1505:note_<=20'b11001100000000000000;
1506:note_<=20'b00101000001111111011;
1507:note_<=20'b01001100000000000000;
1508:note_<=20'b10100100011111101010;
1509:note_<=20'b11000100000000000000;
1510:note_<=20'b00100100010000011010;
1511:note_<=20'b01000100000000000000;
1512:note_<=20'b11010110001111111101;
1513:note_<=20'b11100000000000000000;
1514:note_<=20'b01010100001111110011;
1515:note_<=20'b01100000000000000000;
1516:note_<=20'b11010000000000000001;
1517:note_<=20'b11011100000000000000;
1518:note_<=20'b01010000001111110100;
1519:note_<=20'b01011100000000000000;
1520:note_<=20'b11001100000000000001;
1521:note_<=20'b11011000000000000000;
1522:note_<=20'b01001100010000011010;
1523:note_<=20'b01011000000000000000;
1524:note_<=20'b11000000000000000001;
1525:note_<=20'b11010000000000000000;
1526:note_<=20'b01000000001111111011;
1527:note_<=20'b01010000000000000000;
1528:note_<=20'b11000100001111110101;
1529:note_<=20'b11010100000000000000;
1530:note_<=20'b01000100001111110100;
1531:note_<=20'b01010100000000000000;
1532:note_<=20'b10100100010000011100;
1533:note_<=20'b10110100000000000000;
1534:note_<=20'b00100100001111111011;
1535:note_<=20'b00110100000000000000;
1536:note_<=20'b10101000000000000001;
1537:note_<=20'b10111000000000000000;
1538:note_<=20'b00101000001111110011;
1539:note_<=20'b00111000000000000000;
1540:note_<=20'b10110000000000000001;
1541:note_<=20'b11000100000000000000;
1542:note_<=20'b00110000001111110100;
1543:note_<=20'b01000100000000000000;
1544:note_<=20'b10010100010000011100;
1545:note_<=20'b10111000000000000000;
1546:note_<=20'b00010100001111111011;
1547:note_<=20'b00111000000000000000;
1548:note_<=20'b10100100000000000001;
1549:note_<=20'b11000100000000000000;
1550:note_<=20'b00100100001111110011;
1551:note_<=20'b01000100000000000000;
1552:note_<=20'b10101000000000000001;
1553:note_<=20'b11001100000000000000;
1554:note_<=20'b00101000001111110100;
1555:note_<=20'b01001100000000000000;
1556:note_<=20'b11010100100000011000;
1557:note_<=20'b11100000000000000000;
1558:note_<=20'b01010100001111110011;
1559:note_<=20'b01100000000000000000;
1560:note_<=20'b11010000000000000001;
1561:note_<=20'b11011100000000000000;
1562:note_<=20'b01010000001111110100;
1563:note_<=20'b01011100000000000000;
1564:note_<=20'b11001100000000000001;
1565:note_<=20'b11011000000000000000;
1566:note_<=20'b01001100010000011010;
1567:note_<=20'b01011000000000000000;
1568:note_<=20'b11000000000000000001;
1569:note_<=20'b11010000000000000000;
1570:note_<=20'b01000000001111111011;
1571:note_<=20'b01010000000000000000;
1572:note_<=20'b11000100001111110101;
1573:note_<=20'b11010100000000000000;
1574:note_<=20'b01000100001111110100;
1575:note_<=20'b01010100000000000000;
1576:note_<=20'b11011000010000011100;
1577:note_<=20'b11100000000000000000;
1578:note_<=20'b11110100000000000000;
1579:note_<=20'b01011000001111111011;
1580:note_<=20'b01100000000000000000;
1581:note_<=20'b01110100000000000000;
1582:note_<=20'b11011000001111110101;
1583:note_<=20'b11100000000000000000;
1584:note_<=20'b11110100000000000000;
1585:note_<=20'b01011000001111110100;
1586:note_<=20'b01100000000000000000;
1587:note_<=20'b01110100000000000000;
1588:note_<=20'b11011000000000000001;
1589:note_<=20'b11100000000000000000;
1590:note_<=20'b11110100000000000000;
1591:note_<=20'b01011000010000011010;
1592:note_<=20'b01100000000000000000;
1593:note_<=20'b01110100000000000000;
1594:note_<=20'b11010101001111111101;
1595:note_<=20'b11100000000000000000;
1596:note_<=20'b01010100001111110011;
1597:note_<=20'b01100000000000000000;
1598:note_<=20'b11010000000000000001;
1599:note_<=20'b11011100000000000000;
1600:note_<=20'b01010000001111110100;
1601:note_<=20'b01011100000000000000;
1602:note_<=20'b11001100000000000001;
1603:note_<=20'b11011000000000000000;
1604:note_<=20'b01001100010000011010;
1605:note_<=20'b01011000000000000000;
1606:note_<=20'b11000000000000000001;
1607:note_<=20'b11010000000000000000;
1608:note_<=20'b01000000001111111011;
1609:note_<=20'b01010000000000000000;
1610:note_<=20'b11000100001111110101;
1611:note_<=20'b11010100000000000000;
1612:note_<=20'b01000100001111110100;
1613:note_<=20'b01010100000000000000;
1614:note_<=20'b10100100010000011100;
1615:note_<=20'b10110100000000000000;
1616:note_<=20'b00100100001111111011;
1617:note_<=20'b00110100000000000000;
1618:note_<=20'b10101000000000000001;
1619:note_<=20'b10111000000000000000;
1620:note_<=20'b00101000001111110011;
1621:note_<=20'b00111000000000000000;
1622:note_<=20'b10110000000000000001;
1623:note_<=20'b11000100000000000000;
1624:note_<=20'b00110000001111110100;
1625:note_<=20'b01000100000000000000;
1626:note_<=20'b10010100010000011100;
1627:note_<=20'b10111000000000000000;
1628:note_<=20'b00010100001111111011;
1629:note_<=20'b00111000000000000000;
1630:note_<=20'b10100100000000000001;
1631:note_<=20'b11000100000000000000;
1632:note_<=20'b00100100001111110011;
1633:note_<=20'b01000100000000000000;
1634:note_<=20'b10101000000000000001;
1635:note_<=20'b11001100000000000000;
1636:note_<=20'b00101000001111110100;
1637:note_<=20'b01001100000000000000;
1638:note_<=20'b10110100100000011000;
1639:note_<=20'b11010000000000000000;
1640:note_<=20'b00110100001111110011;
1641:note_<=20'b01010000000000000000;
1642:note_<=20'b10101000100000010001;
1643:note_<=20'b11001100000000000000;
1644:note_<=20'b00101000001111111011;
1645:note_<=20'b01001100000000000000;
1646:note_<=20'b10100100011111101010;
1647:note_<=20'b11000100000000000000;
1648:note_<=20'b00100100010000011010;
1649:note_<=20'b01000100000000000000;
1650:note_<=20'b10110101101111100110;
1651:note_<=20'b11000100000000000000;
1652:note_<=20'b00110100010000011010;
1653:note_<=20'b01000100000000000000;
1654:note_<=20'b10110100000000000001;
1655:note_<=20'b11000100000000000000;
1656:note_<=20'b00110100001111111011;
1657:note_<=20'b01000100000000000000;
1658:note_<=20'b10110100001111110101;
1659:note_<=20'b11000100000000000000;
1660:note_<=20'b00110100001111110100;
1661:note_<=20'b01000100000000000000;
1662:note_<=20'b10110100010000011100;
1663:note_<=20'b11000100000000000000;
1664:note_<=20'b00110100001111111011;
1665:note_<=20'b01000100000000000000;
1666:note_<=20'b10111100000000000001;
1667:note_<=20'b11001100000000000000;
1668:note_<=20'b00111100001111110011;
1669:note_<=20'b01001100000000000000;
1670:note_<=20'b10110000001111110110;
1671:note_<=20'b11010100000000000000;
1672:note_<=20'b00110000010000011010;
1673:note_<=20'b01010100000000000000;
1674:note_<=20'b10100100000000000001;
1675:note_<=20'b11000100000000000000;
1676:note_<=20'b00100100001111111011;
1677:note_<=20'b01000100000000000000;
1678:note_<=20'b10100100001111110101;
1679:note_<=20'b10111000000000000000;
1680:note_<=20'b00100100001111110100;
1681:note_<=20'b00111000000000000000;
1682:note_<=20'b10010100000000000001;
1683:note_<=20'b10110000000000000000;
1684:note_<=20'b00010100010000011010;
1685:note_<=20'b00110000000000000000;
1686:note_<=20'b10110100101111100110;
1687:note_<=20'b11000100000000000000;
1688:note_<=20'b00110100010000011010;
1689:note_<=20'b01000100000000000000;
1690:note_<=20'b10110100000000000001;
1691:note_<=20'b11000100000000000000;
1692:note_<=20'b00110100001111111011;
1693:note_<=20'b01000100000000000000;
1694:note_<=20'b10110100001111110101;
1695:note_<=20'b11000100000000000000;
1696:note_<=20'b00110100001111110100;
1697:note_<=20'b01000100000000000000;
1698:note_<=20'b10110100010000011100;
1699:note_<=20'b11000100000000000000;
1700:note_<=20'b00110100001111111011;
1701:note_<=20'b01000100000000000000;
1702:note_<=20'b10111100000000000001;
1703:note_<=20'b11001100000000000000;
1704:note_<=20'b00111100001111110011;
1705:note_<=20'b01001100000000000000;
1706:note_<=20'b10110000000000000001;
1707:note_<=20'b11010100000000000000;
1708:note_<=20'b00110000001111110100;
1709:note_<=20'b01010100000000000000;
1710:note_<=20'b10110110000000000001;
1711:note_<=20'b11000100000000000000;
1712:note_<=20'b00110100010000011010;
1713:note_<=20'b01000100000000000000;
1714:note_<=20'b10110100000000000001;
1715:note_<=20'b11000100000000000000;
1716:note_<=20'b00110100001111111011;
1717:note_<=20'b01000100000000000000;
1718:note_<=20'b10110100001111110101;
1719:note_<=20'b11000100000000000000;
1720:note_<=20'b00110100001111110100;
1721:note_<=20'b01000100000000000000;
1722:note_<=20'b10110100010000011100;
1723:note_<=20'b11000100000000000000;
1724:note_<=20'b00110100001111111011;
1725:note_<=20'b01000100000000000000;
1726:note_<=20'b10111100000000000001;
1727:note_<=20'b11001100000000000000;
1728:note_<=20'b00111100001111110011;
1729:note_<=20'b01001100000000000000;
1730:note_<=20'b10110000001111110110;
1731:note_<=20'b11010100000000000000;
1732:note_<=20'b00110000010000011010;
1733:note_<=20'b01010100000000000000;
1734:note_<=20'b10100100000000000001;
1735:note_<=20'b11000100000000000000;
1736:note_<=20'b00100100001111111011;
1737:note_<=20'b01000100000000000000;
1738:note_<=20'b10100100001111110101;
1739:note_<=20'b10111000000000000000;
1740:note_<=20'b00100100001111110100;
1741:note_<=20'b00111000000000000000;
1742:note_<=20'b10010100000000000001;
1743:note_<=20'b10110000000000000000;
1744:note_<=20'b00010100010000011010;
1745:note_<=20'b00110000000000000000;
1746:note_<=20'b10101100101111100110;
1747:note_<=20'b11010100000000000000;
1748:note_<=20'b00101100010000011010;
1749:note_<=20'b01010100000000000000;
1750:note_<=20'b10101100000000000001;
1751:note_<=20'b11010100000000000000;
1752:note_<=20'b00101100001111111011;
1753:note_<=20'b01010100000000000000;
1754:note_<=20'b10101100001111110101;
1755:note_<=20'b11010100000000000000;
1756:note_<=20'b00101100001111110100;
1757:note_<=20'b01010100000000000000;
1758:note_<=20'b10101100010000011100;
1759:note_<=20'b11000100000000000000;
1760:note_<=20'b00101100001111111011;
1761:note_<=20'b01000100000000000000;
1762:note_<=20'b10101100000000000001;
1763:note_<=20'b11010100000000000000;
1764:note_<=20'b00101100001111110011;
1765:note_<=20'b01010100000000000000;
1766:note_<=20'b10110000001111110110;
1767:note_<=20'b11000000000000000000;
1768:note_<=20'b11100000000000000000;
1769:note_<=20'b00110000010000011010;
1770:note_<=20'b01000000000000000000;
1771:note_<=20'b01100000000000000000;
1772:note_<=20'b10110000101111100110;
1773:note_<=20'b00110000010000011010;
1774:note_<=20'b10100100101111100110;
1775:note_<=20'b11000100000000000000;
1776:note_<=20'b00100100010000011010;
1777:note_<=20'b01000100000000000000;
1778:note_<=20'b10010100011111110001;
1779:note_<=20'b10110000000000000000;
1780:note_<=20'b00010100001111110100;
1781:note_<=20'b00110000000000000000;
1782:note_<=20'b10000000100000011000;
1783:note_<=20'b10100100000000000000;
1784:note_<=20'b00000000001111110011;
1785:note_<=20'b00100100000000000000;
1786:note_<=20'b10010100100000010001;
1787:note_<=20'b10111000000000000000;
1788:note_<=20'b00010100001111111011;
1789:note_<=20'b00111000000000000000;
1790:note_<=20'b10011100001111110101;
1791:note_<=20'b11000000000000000000;
1792:note_<=20'b00011100001111110100;
1793:note_<=20'b01000000000000000000;
1794:note_<=20'b10011000010000011100;
1795:note_<=20'b10111100000000000000;
1796:note_<=20'b00011000001111111011;
1797:note_<=20'b00111100000000000000;
1798:note_<=20'b10010100000000000001;
1799:note_<=20'b10111000000000000000;
1800:note_<=20'b00010100001111110011;
1801:note_<=20'b00111000000000000000;
1802:note_<=20'b10010100001111110110;
1803:note_<=20'b10110000000000000000;
1804:note_<=20'b00010100001011000000;
1805:note_<=20'b00110000000000000000;
1806:note_<=20'b10110000001010101011;
1807:note_<=20'b11010100000000000000;
1808:note_<=20'b00110000001010101001;
1809:note_<=20'b01010100000000000000;
1810:note_<=20'b11000000001010101100;
1811:note_<=20'b11100000000000000000;
1812:note_<=20'b01000000001010010101;
1813:note_<=20'b01100000000000000000;
1814:note_<=20'b11000100001010101011;
1815:note_<=20'b11101000000000000000;
1816:note_<=20'b01000100010000011010;
1817:note_<=20'b01101000000000000000;
1818:note_<=20'b10111000001111111101;
1819:note_<=20'b11011000000000000000;
1820:note_<=20'b00111000001111110011;
1821:note_<=20'b01011000000000000000;
1822:note_<=20'b11000000000000000001;
1823:note_<=20'b11100000000000000000;
1824:note_<=20'b01000000001111110100;
1825:note_<=20'b01100000000000000000;
1826:note_<=20'b10111000010000011100;
1827:note_<=20'b11010100000000000000;
1828:note_<=20'b00111000001111111011;
1829:note_<=20'b01010100000000000000;
1830:note_<=20'b10100100001111110101;
1831:note_<=20'b11000100000000000000;
1832:note_<=20'b00100100001111110100;
1833:note_<=20'b01000100000000000000;
1834:note_<=20'b10101000000000000001;
1835:note_<=20'b11001100000000000000;
1836:note_<=20'b00101000010000011010;
1837:note_<=20'b01001100000000000000;
1838:note_<=20'b10011100000000000001;
1839:note_<=20'b11000000000000000000;
1840:note_<=20'b00011100001111111011;
1841:note_<=20'b01000000000000000000;
1842:note_<=20'b10100100011111101010;
1843:note_<=20'b11000100000000000000;
1844:note_<=20'b00100100010000011010;
1845:note_<=20'b01000100000000000000;
1846:note_<=20'b10010100011111110001;
1847:note_<=20'b10110000000000000000;
1848:note_<=20'b00010100001111110100;
1849:note_<=20'b00110000000000000000;
1850:note_<=20'b10000000100000011000;
1851:note_<=20'b10100100000000000000;
1852:note_<=20'b00000000001111110011;
1853:note_<=20'b00100100000000000000;
1854:note_<=20'b10010100100000010001;
1855:note_<=20'b10111000000000000000;
1856:note_<=20'b00010100001111111011;
1857:note_<=20'b00111000000000000000;
1858:note_<=20'b10011100001111110101;
1859:note_<=20'b11000000000000000000;
1860:note_<=20'b00011100001111110100;
1861:note_<=20'b01000000000000000000;
1862:note_<=20'b10011000010000011100;
1863:note_<=20'b10111100000000000000;
1864:note_<=20'b00011000001111111011;
1865:note_<=20'b00111100000000000000;
1866:note_<=20'b10010100000000000001;
1867:note_<=20'b10111000000000000000;
1868:note_<=20'b00010100001111110011;
1869:note_<=20'b00111000000000000000;
1870:note_<=20'b10010100001111110110;
1871:note_<=20'b10110000000000000000;
1872:note_<=20'b00010100001011000000;
1873:note_<=20'b00110000000000000000;
1874:note_<=20'b10110000001010101011;
1875:note_<=20'b11010100000000000000;
1876:note_<=20'b00110000001010101001;
1877:note_<=20'b01010100000000000000;
1878:note_<=20'b11000000001010101100;
1879:note_<=20'b11100000000000000000;
1880:note_<=20'b01000000001010010101;
1881:note_<=20'b01100000000000000000;
1882:note_<=20'b11000100001010101011;
1883:note_<=20'b11101000000000000000;
1884:note_<=20'b01000100010000011010;
1885:note_<=20'b01101000000000000000;
1886:note_<=20'b10111000001111111101;
1887:note_<=20'b11011000000000000000;
1888:note_<=20'b00111000001111110011;
1889:note_<=20'b01011000000000000000;
1890:note_<=20'b11000000000000000001;
1891:note_<=20'b11100000000000000000;
1892:note_<=20'b01000000001111110100;
1893:note_<=20'b01100000000000000000;
1894:note_<=20'b10111000010000011100;
1895:note_<=20'b11010100000000000000;
1896:note_<=20'b00111000001111111011;
1897:note_<=20'b01010100000000000000;
1898:note_<=20'b10100100001111110101;
1899:note_<=20'b11000100000000000000;
1900:note_<=20'b00100100001111110100;
1901:note_<=20'b01000100000000000000;
1902:note_<=20'b10101000000000000001;
1903:note_<=20'b11001100000000000000;
1904:note_<=20'b00101000010000011010;
1905:note_<=20'b01001100000000000000;
1906:note_<=20'b10011100000000000001;
1907:note_<=20'b11000000000000000000;
1908:note_<=20'b00011100001111111011;
1909:note_<=20'b01000000000000000000;
1910:note_<=20'b11000100011111101010;
1911:note_<=20'b11010100000000000000;
1912:note_<=20'b01000100010000011010;
1913:note_<=20'b01010100000000000000;
1914:note_<=20'b10111000000000000001;
1915:note_<=20'b11000100000000000000;
1916:note_<=20'b00111000001111111011;
1917:note_<=20'b01000100000000000000;
1918:note_<=20'b10100100001111110101;
1919:note_<=20'b10110000000000000000;
1920:note_<=20'b00100100001111110100;
1921:note_<=20'b00110000000000000000;
1922:note_<=20'b10100100100000011000;
1923:note_<=20'b10110100000000000000;
1924:note_<=20'b00100100001111110011;
1925:note_<=20'b00110100000000000000;
1926:note_<=20'b10101000001111110110;
1927:note_<=20'b10111000000000000000;
1928:note_<=20'b00101000010000011010;
1929:note_<=20'b00111000000000000000;
1930:note_<=20'b11000100000000000001;
1931:note_<=20'b11011000000000000000;
1932:note_<=20'b01000100001111111011;
1933:note_<=20'b01011000000000000000;
1934:note_<=20'b11000100001111110101;
1935:note_<=20'b11011000000000000000;
1936:note_<=20'b01000100001111110100;
1937:note_<=20'b01011000000000000000;
1938:note_<=20'b10101000000000000001;
1939:note_<=20'b10111000000000000000;
1940:note_<=20'b00101000010000011010;
1941:note_<=20'b00111000000000000000;
1942:note_<=20'b10110000101111100110;
1943:note_<=20'b11000000000000000000;
1944:note_<=20'b00110000001011000000;
1945:note_<=20'b01000000000000000000;
1946:note_<=20'b11011000001010101011;
1947:note_<=20'b11101000000000000000;
1948:note_<=20'b01011000001010101001;
1949:note_<=20'b01101000000000000000;
1950:note_<=20'b11011000001010101100;
1951:note_<=20'b11101000000000000000;
1952:note_<=20'b01011000001010010101;
1953:note_<=20'b01101000000000000000;
1954:note_<=20'b11011000001010101011;
1955:note_<=20'b11101000000000000000;
1956:note_<=20'b01011000001011000000;
1957:note_<=20'b01101000000000000000;
1958:note_<=20'b11010100001010101011;
1959:note_<=20'b11100000000000000000;
1960:note_<=20'b01010100001010101001;
1961:note_<=20'b01100000000000000000;
1962:note_<=20'b11001100001010101100;
1963:note_<=20'b11011000000000000000;
1964:note_<=20'b01001100001010010101;
1965:note_<=20'b01011000000000000000;
1966:note_<=20'b11000100001010101011;
1967:note_<=20'b11010100000000000000;
1968:note_<=20'b01000100010000011010;
1969:note_<=20'b01010100000000000000;
1970:note_<=20'b10111000000000000001;
1971:note_<=20'b11000100000000000000;
1972:note_<=20'b00111000001111111011;
1973:note_<=20'b01000100000000000000;
1974:note_<=20'b10101000001111110101;
1975:note_<=20'b10111000000000000000;
1976:note_<=20'b00101000001111110100;
1977:note_<=20'b00111000000000000000;
1978:note_<=20'b10100100000000000001;
1979:note_<=20'b10110000000000000000;
1980:note_<=20'b00100100010000011010;
1981:note_<=20'b00110000000000000000;
1982:note_<=20'b11000100101111100110;
1983:note_<=20'b11010100000000000000;
1984:note_<=20'b01000100010000011010;
1985:note_<=20'b01010100000000000000;
1986:note_<=20'b10111000000000000001;
1987:note_<=20'b11000100000000000000;
1988:note_<=20'b00111000001111111011;
1989:note_<=20'b01000100000000000000;
1990:note_<=20'b10100100001111110101;
1991:note_<=20'b10110000000000000000;
1992:note_<=20'b00100100001111110100;
1993:note_<=20'b00110000000000000000;
1994:note_<=20'b10100100100000011000;
1995:note_<=20'b10110100000000000000;
1996:note_<=20'b00100100001111110011;
1997:note_<=20'b00110100000000000000;
1998:note_<=20'b10101000001111110110;
1999:note_<=20'b10111000000000000000;
2000:note_<=20'b00101000010000011010;
2001:note_<=20'b00111000000000000000;
2002:note_<=20'b11000100000000000001;
2003:note_<=20'b11011000000000000000;
2004:note_<=20'b01000100001111111011;
2005:note_<=20'b01011000000000000000;
2006:note_<=20'b11000100001111110101;
2007:note_<=20'b11011000000000000000;
2008:note_<=20'b01000100001111110100;
2009:note_<=20'b01011000000000000000;
2010:note_<=20'b10101000000000000001;
2011:note_<=20'b10111000000000000000;
2012:note_<=20'b00101000010000011010;
2013:note_<=20'b00111000000000000000;
2014:note_<=20'b10110000101111100110;
2015:note_<=20'b11000000000000000000;
2016:note_<=20'b00110000010000011010;
2017:note_<=20'b01000000000000000000;
2018:note_<=20'b11001100000000000001;
2019:note_<=20'b11011000000000000000;
2020:note_<=20'b01001100001111111011;
2021:note_<=20'b01011000000000000000;
2022:note_<=20'b11001100001111110101;
2023:note_<=20'b11011000000000000000;
2024:note_<=20'b01001100001111110100;
2025:note_<=20'b01011000000000000000;
2026:note_<=20'b11001100000000000001;
2027:note_<=20'b11011000000000000000;
2028:note_<=20'b01001100001011000000;
2029:note_<=20'b01011000000000000000;
2030:note_<=20'b11000100001010101011;
2031:note_<=20'b11010100000000000000;
2032:note_<=20'b01000100001010101001;
2033:note_<=20'b01010100000000000000;
2034:note_<=20'b11000000001010101100;
2035:note_<=20'b11001100000000000000;
2036:note_<=20'b01000000001010010101;
2037:note_<=20'b01001100000000000000;
2038:note_<=20'b10110000001010101011;
2039:note_<=20'b11000100000000000000;
2040:note_<=20'b00110000010000011010;
2041:note_<=20'b01000100000000000000;
2042:note_<=20'b10100100000000000001;
2043:note_<=20'b00100100001111111011;
2044:note_<=20'b10100100001111110101;
2045:note_<=20'b00100100001111110100;
2046:note_<=20'b10010100000000000001;
2047:note_<=20'b00010100010000011010;
2048:note_<=20'b11000100101111100110;
2049:note_<=20'b11010100000000000000;
2050:note_<=20'b01000100010000011010;
2051:note_<=20'b01010100000000000000;
2052:note_<=20'b10111000000000000001;
2053:note_<=20'b11000100000000000000;
2054:note_<=20'b00111000001111111011;
2055:note_<=20'b01000100000000000000;
2056:note_<=20'b10100100001111110101;
2057:note_<=20'b10110000000000000000;
2058:note_<=20'b00100100001111110100;
2059:note_<=20'b00110000000000000000;
2060:note_<=20'b10100100100000011000;
2061:note_<=20'b10110100000000000000;
2062:note_<=20'b00100100001111110011;
2063:note_<=20'b00110100000000000000;
2064:note_<=20'b10101000001111110110;
2065:note_<=20'b10111000000000000000;
2066:note_<=20'b00101000010000011010;
2067:note_<=20'b00111000000000000000;
2068:note_<=20'b11000100000000000001;
2069:note_<=20'b11011000000000000000;
2070:note_<=20'b01000100001111111011;
2071:note_<=20'b01011000000000000000;
2072:note_<=20'b11000100001111110101;
2073:note_<=20'b11011000000000000000;
2074:note_<=20'b01000100001111110100;
2075:note_<=20'b01011000000000000000;
2076:note_<=20'b10101000000000000001;
2077:note_<=20'b10111000000000000000;
2078:note_<=20'b00101000010000011010;
2079:note_<=20'b00111000000000000000;
2080:note_<=20'b10110000101111100110;
2081:note_<=20'b11000000000000000000;
2082:note_<=20'b00110000001011000000;
2083:note_<=20'b01000000000000000000;
2084:note_<=20'b11011000001010101011;
2085:note_<=20'b11101000000000000000;
2086:note_<=20'b01011000001010101001;
2087:note_<=20'b01101000000000000000;
2088:note_<=20'b11011000001010101100;
2089:note_<=20'b11101000000000000000;
2090:note_<=20'b01011000001010010101;
2091:note_<=20'b01101000000000000000;
2092:note_<=20'b11011000001010101011;
2093:note_<=20'b11101000000000000000;
2094:note_<=20'b01011000001011000000;
2095:note_<=20'b01101000000000000000;
2096:note_<=20'b11010100001010101011;
2097:note_<=20'b11100000000000000000;
2098:note_<=20'b01010100001010101001;
2099:note_<=20'b01100000000000000000;
2100:note_<=20'b11001100001010101100;
2101:note_<=20'b11011000000000000000;
2102:note_<=20'b01001100001010010101;
2103:note_<=20'b01011000000000000000;
2104:note_<=20'b11000100001010101011;
2105:note_<=20'b11010100000000000000;
2106:note_<=20'b01000100010000011010;
2107:note_<=20'b01010100000000000000;
2108:note_<=20'b10111000000000000001;
2109:note_<=20'b11000100000000000000;
2110:note_<=20'b00111000001111111011;
2111:note_<=20'b01000100000000000000;
2112:note_<=20'b10101000001111110101;
2113:note_<=20'b10111000000000000000;
2114:note_<=20'b00101000001111110100;
2115:note_<=20'b00111000000000000000;
2116:note_<=20'b10100100000000000001;
2117:note_<=20'b10110000000000000000;
2118:note_<=20'b00100100010000011010;
2119:note_<=20'b00110000000000000000;
2120:note_<=20'b11000100101111100110;
2121:note_<=20'b11010100000000000000;
2122:note_<=20'b01000100010000011010;
2123:note_<=20'b01010100000000000000;
2124:note_<=20'b10111000000000000001;
2125:note_<=20'b11000100000000000000;
2126:note_<=20'b00111000001111111011;
2127:note_<=20'b01000100000000000000;
2128:note_<=20'b10100100001111110101;
2129:note_<=20'b10110000000000000000;
2130:note_<=20'b00100100001111110100;
2131:note_<=20'b00110000000000000000;
2132:note_<=20'b10100100100000011000;
2133:note_<=20'b10110100000000000000;
2134:note_<=20'b00100100001111110011;
2135:note_<=20'b00110100000000000000;
2136:note_<=20'b10101000001111110110;
2137:note_<=20'b10111000000000000000;
2138:note_<=20'b00101000010000011010;
2139:note_<=20'b00111000000000000000;
2140:note_<=20'b11000100000000000001;
2141:note_<=20'b11011000000000000000;
2142:note_<=20'b01000100001111111011;
2143:note_<=20'b01011000000000000000;
2144:note_<=20'b11000100001111110101;
2145:note_<=20'b11011000000000000000;
2146:note_<=20'b01000100001111110100;
2147:note_<=20'b01011000000000000000;
2148:note_<=20'b10101000000000000001;
2149:note_<=20'b10111000000000000000;
2150:note_<=20'b00101000010000011010;
2151:note_<=20'b00111000000000000000;
2152:note_<=20'b10110000101111100110;
2153:note_<=20'b11000000000000000000;
2154:note_<=20'b00110000010000011010;
2155:note_<=20'b01000000000000000000;
2156:note_<=20'b11001100000000000001;
2157:note_<=20'b11011000000000000000;
2158:note_<=20'b01001100001111111011;
2159:note_<=20'b01011000000000000000;
2160:note_<=20'b11001100001111110101;
2161:note_<=20'b11011000000000000000;
2162:note_<=20'b01001100001111110100;
2163:note_<=20'b01011000000000000000;
2164:note_<=20'b11001100000000000001;
2165:note_<=20'b11011000000000000000;
2166:note_<=20'b01001100001011000000;
2167:note_<=20'b01011000000000000000;
2168:note_<=20'b11000100001010101011;
2169:note_<=20'b11010100000000000000;
2170:note_<=20'b01000100001010101001;
2171:note_<=20'b01010100000000000000;
2172:note_<=20'b11000000001010101100;
2173:note_<=20'b11001100000000000000;
2174:note_<=20'b01000000001010010101;
2175:note_<=20'b01001100000000000000;
2176:note_<=20'b10110000001010101011;
2177:note_<=20'b11000100000000000000;
2178:note_<=20'b00110000010000011010;
2179:note_<=20'b01000100000000000000;
2180:note_<=20'b10100100000000000001;
2181:note_<=20'b00100100001111111011;
2182:note_<=20'b10100100001111110101;
2183:note_<=20'b00100100001111110100;
2184:note_<=20'b10010100000000000001;
2185:note_<=20'b00010100010000011010;
2186:note_<=20'b10110100101111100110;
2187:note_<=20'b11000100000000000000;
2188:note_<=20'b00110100010000011010;
2189:note_<=20'b01000100000000000000;
2190:note_<=20'b10110100000000000001;
2191:note_<=20'b11000100000000000000;
2192:note_<=20'b00110100001111111011;
2193:note_<=20'b01000100000000000000;
2194:note_<=20'b10110100001111110101;
2195:note_<=20'b11000100000000000000;
2196:note_<=20'b00110100001111110100;
2197:note_<=20'b01000100000000000000;
2198:note_<=20'b10110100010000011100;
2199:note_<=20'b11000100000000000000;
2200:note_<=20'b00110100001111111011;
2201:note_<=20'b01000100000000000000;
2202:note_<=20'b10111100000000000001;
2203:note_<=20'b11001100000000000000;
2204:note_<=20'b00111100001111110011;
2205:note_<=20'b01001100000000000000;
2206:note_<=20'b10110000001111110110;
2207:note_<=20'b11010100000000000000;
2208:note_<=20'b00110000010000011010;
2209:note_<=20'b01010100000000000000;
2210:note_<=20'b10100100000000000001;
2211:note_<=20'b11000100000000000000;
2212:note_<=20'b00100100001111111011;
2213:note_<=20'b01000100000000000000;
2214:note_<=20'b10100100001111110101;
2215:note_<=20'b10111000000000000000;
2216:note_<=20'b00100100001111110100;
2217:note_<=20'b00111000000000000000;
2218:note_<=20'b10010100000000000001;
2219:note_<=20'b10110000000000000000;
2220:note_<=20'b00010100010000011010;
2221:note_<=20'b00110000000000000000;
2222:note_<=20'b10110100101111100110;
2223:note_<=20'b11000100000000000000;
2224:note_<=20'b00110100010000011010;
2225:note_<=20'b01000100000000000000;
2226:note_<=20'b10110100000000000001;
2227:note_<=20'b11000100000000000000;
2228:note_<=20'b00110100001111111011;
2229:note_<=20'b01000100000000000000;
2230:note_<=20'b10110100001111110101;
2231:note_<=20'b11000100000000000000;
2232:note_<=20'b00110100001111110100;
2233:note_<=20'b01000100000000000000;
2234:note_<=20'b10110100010000011100;
2235:note_<=20'b11000100000000000000;
2236:note_<=20'b00110100001111111011;
2237:note_<=20'b01000100000000000000;
2238:note_<=20'b10111100000000000001;
2239:note_<=20'b11001100000000000000;
2240:note_<=20'b00111100001111110011;
2241:note_<=20'b01001100000000000000;
2242:note_<=20'b10110000000000000001;
2243:note_<=20'b11010100000000000000;
2244:note_<=20'b00110000001111110100;
2245:note_<=20'b01010100000000000000;
2246:note_<=20'b10110110000000000001;
2247:note_<=20'b11000100000000000000;
2248:note_<=20'b00110100010000011010;
2249:note_<=20'b01000100000000000000;
2250:note_<=20'b10110100000000000001;
2251:note_<=20'b11000100000000000000;
2252:note_<=20'b00110100001111111011;
2253:note_<=20'b01000100000000000000;
2254:note_<=20'b10110100001111110101;
2255:note_<=20'b11000100000000000000;
2256:note_<=20'b00110100001111110100;
2257:note_<=20'b01000100000000000000;
2258:note_<=20'b10110100010000011100;
2259:note_<=20'b11000100000000000000;
2260:note_<=20'b00110100001111111011;
2261:note_<=20'b01000100000000000000;
2262:note_<=20'b10111100000000000001;
2263:note_<=20'b11001100000000000000;
2264:note_<=20'b00111100001111110011;
2265:note_<=20'b01001100000000000000;
2266:note_<=20'b10110000001111110110;
2267:note_<=20'b11010100000000000000;
2268:note_<=20'b00110000010000011010;
2269:note_<=20'b01010100000000000000;
2270:note_<=20'b10100100000000000001;
2271:note_<=20'b11000100000000000000;
2272:note_<=20'b00100100001111111011;
2273:note_<=20'b01000100000000000000;
2274:note_<=20'b10100100001111110101;
2275:note_<=20'b10111000000000000000;
2276:note_<=20'b00100100001111110100;
2277:note_<=20'b00111000000000000000;
2278:note_<=20'b10010100000000000001;
2279:note_<=20'b10110000000000000000;
2280:note_<=20'b00010100010000011010;
2281:note_<=20'b00110000000000000000;
2282:note_<=20'b10101100101111100110;
2283:note_<=20'b11010100000000000000;
2284:note_<=20'b00101100010000011010;
2285:note_<=20'b01010100000000000000;
2286:note_<=20'b10101100000000000001;
2287:note_<=20'b11010100000000000000;
2288:note_<=20'b00101100001111111011;
2289:note_<=20'b01010100000000000000;
2290:note_<=20'b10101100001111110101;
2291:note_<=20'b11010100000000000000;
2292:note_<=20'b00101100001111110100;
2293:note_<=20'b01010100000000000000;
2294:note_<=20'b10101100010000011100;
2295:note_<=20'b11000100000000000000;
2296:note_<=20'b00101100001111111011;
2297:note_<=20'b01000100000000000000;
2298:note_<=20'b10101100000000000001;
2299:note_<=20'b11010100000000000000;
2300:note_<=20'b00101100001111110011;
2301:note_<=20'b01010100000000000000;
2302:note_<=20'b10110000001111110110;
2303:note_<=20'b11000000000000000000;
2304:note_<=20'b11100000000000000000;
2305:note_<=20'b00110000010000011010;
2306:note_<=20'b01000000000000000000;
2307:note_<=20'b01100000000000000000;
2308:note_<=20'b10110000101111100110;
2309:note_<=20'b00110000010000011010;
2310:note_<=20'b11000100101111100110;
2311:note_<=20'b11010100000000000000;
2312:note_<=20'b01000100010000011010;
2313:note_<=20'b01010100000000000000;
2314:note_<=20'b10111000000000000001;
2315:note_<=20'b11000100000000000000;
2316:note_<=20'b00111000001111111011;
2317:note_<=20'b01000100000000000000;
2318:note_<=20'b10100100001111110101;
2319:note_<=20'b10110000000000000000;
2320:note_<=20'b00100100001111110100;
2321:note_<=20'b00110000000000000000;
2322:note_<=20'b10100100100000011000;
2323:note_<=20'b10110100000000000000;
2324:note_<=20'b00100100001111110011;
2325:note_<=20'b00110100000000000000;
2326:note_<=20'b10101000001111110110;
2327:note_<=20'b10111000000000000000;
2328:note_<=20'b00101000010000011010;
2329:note_<=20'b00111000000000000000;
2330:note_<=20'b11000100000000000001;
2331:note_<=20'b11011000000000000000;
2332:note_<=20'b01000100001111111011;
2333:note_<=20'b01011000000000000000;
2334:note_<=20'b11000100001111110101;
2335:note_<=20'b11011000000000000000;
2336:note_<=20'b01000100001111110100;
2337:note_<=20'b01011000000000000000;
2338:note_<=20'b10101000000000000001;
2339:note_<=20'b10111000000000000000;
2340:note_<=20'b00101000010000011010;
2341:note_<=20'b00111000000000000000;
2342:note_<=20'b10110000101111100110;
2343:note_<=20'b11000000000000000000;
2344:note_<=20'b00110000001011000000;
2345:note_<=20'b01000000000000000000;
2346:note_<=20'b11011000001010101011;
2347:note_<=20'b11101000000000000000;
2348:note_<=20'b01011000001010101001;
2349:note_<=20'b01101000000000000000;
2350:note_<=20'b11011000001010101100;
2351:note_<=20'b11101000000000000000;
2352:note_<=20'b01011000001010010101;
2353:note_<=20'b01101000000000000000;
2354:note_<=20'b11011000001010101011;
2355:note_<=20'b11101000000000000000;
2356:note_<=20'b01011000001011000000;
2357:note_<=20'b01101000000000000000;
2358:note_<=20'b11010100001010101011;
2359:note_<=20'b11100000000000000000;
2360:note_<=20'b01010100001010101001;
2361:note_<=20'b01100000000000000000;
2362:note_<=20'b11001100001010101100;
2363:note_<=20'b11011000000000000000;
2364:note_<=20'b01001100001010010101;
2365:note_<=20'b01011000000000000000;
2366:note_<=20'b11000100001010101011;
2367:note_<=20'b11010100000000000000;
2368:note_<=20'b01000100010000011010;
2369:note_<=20'b01010100000000000000;
2370:note_<=20'b10111000000000000001;
2371:note_<=20'b11000100000000000000;
2372:note_<=20'b00111000001111111011;
2373:note_<=20'b01000100000000000000;
2374:note_<=20'b10101000001111110101;
2375:note_<=20'b10111000000000000000;
2376:note_<=20'b00101000001111110100;
2377:note_<=20'b00111000000000000000;
2378:note_<=20'b10100100000000000001;
2379:note_<=20'b10110000000000000000;
2380:note_<=20'b00100100010000011010;
2381:note_<=20'b00110000000000000000;
2382:note_<=20'b11000100101111100110;
2383:note_<=20'b11010100000000000000;
2384:note_<=20'b01000100010000011010;
2385:note_<=20'b01010100000000000000;
2386:note_<=20'b10111000000000000001;
2387:note_<=20'b11000100000000000000;
2388:note_<=20'b00111000001111111011;
2389:note_<=20'b01000100000000000000;
2390:note_<=20'b10100100001111110101;
2391:note_<=20'b10110000000000000000;
2392:note_<=20'b00100100001111110100;
2393:note_<=20'b00110000000000000000;
2394:note_<=20'b10100100100000011000;
2395:note_<=20'b10110100000000000000;
2396:note_<=20'b00100100001111110011;
2397:note_<=20'b00110100000000000000;
2398:note_<=20'b10101000001111110110;
2399:note_<=20'b10111000000000000000;
2400:note_<=20'b00101000010000011010;
2401:note_<=20'b00111000000000000000;
2402:note_<=20'b11000100000000000001;
2403:note_<=20'b11011000000000000000;
2404:note_<=20'b01000100001111111011;
2405:note_<=20'b01011000000000000000;
2406:note_<=20'b11000100001111110101;
2407:note_<=20'b11011000000000000000;
2408:note_<=20'b01000100001111110100;
2409:note_<=20'b01011000000000000000;
2410:note_<=20'b10101000000000000001;
2411:note_<=20'b10111000000000000000;
2412:note_<=20'b00101000010000011010;
2413:note_<=20'b00111000000000000000;
2414:note_<=20'b10110000101111100110;
2415:note_<=20'b11000000000000000000;
2416:note_<=20'b00110000010000011010;
2417:note_<=20'b01000000000000000000;
2418:note_<=20'b11001100000000000001;
2419:note_<=20'b11011000000000000000;
2420:note_<=20'b01001100001111111011;
2421:note_<=20'b01011000000000000000;
2422:note_<=20'b11001100001111110101;
2423:note_<=20'b11011000000000000000;
2424:note_<=20'b01001100001111110100;
2425:note_<=20'b01011000000000000000;
2426:note_<=20'b11001100000000000001;
2427:note_<=20'b11011000000000000000;
2428:note_<=20'b01001100001011000000;
2429:note_<=20'b01011000000000000000;
2430:note_<=20'b11000100001010101011;
2431:note_<=20'b11010100000000000000;
2432:note_<=20'b01000100001010101001;
2433:note_<=20'b01010100000000000000;
2434:note_<=20'b11000000001010101100;
2435:note_<=20'b11001100000000000000;
2436:note_<=20'b01000000001010010101;
2437:note_<=20'b01001100000000000000;
2438:note_<=20'b10110000001010101011;
2439:note_<=20'b11000100000000000000;
2440:note_<=20'b00110000010000011010;
2441:note_<=20'b01000100000000000000;
2442:note_<=20'b10100100000000000001;
2443:note_<=20'b00100100001111111011;
2444:note_<=20'b10100100001111110101;
2445:note_<=20'b00100100001111110100;
2446:note_<=20'b10010100000000000001;
2447:note_<=20'b00010100010000011010;
default: note_ <= 20'b0;
endcase

note_on <= note_[19:19];
note <= note_[18:14];
delay <= note_[13:0];
end
endmodule


